`timescale 1ns/1ns

module wt_fc1_mem7 #(parameter ADDR_WIDTH = 11, DATA_WIDTH = 144, DEPTH = 1024) (
input wire clk,
input wire [ADDR_WIDTH-1:0] addr_a, 
input wire [ADDR_WIDTH-1:0] addr_b, 
output reg [DATA_WIDTH-1:0] q_a,
output reg [DATA_WIDTH-1:0] q_b
);

reg [DATA_WIDTH-1:0] mem [0:DEPTH-1];

initial begin
mem[0] = 144'h00b300aa03d004fb038effeb006f0005038a;
mem[1] = 144'hff440276022affcb00faff24fe8cfd890045;
mem[2] = 144'hfe6b039600aafe61001500f4fe17fd14fe8d;
mem[3] = 144'hff26ff07fcaf023302defd72fcaa01eafe94;
mem[4] = 144'h015d030b02630228037a0143fcfbfe610148;
mem[5] = 144'hfebaff7b00cd017cff43fd95fe0bffc7fe92;
mem[6] = 144'hff3c00de021203c900deffa7fdd6012502c0;
mem[7] = 144'h019eff360169032801060173ffd100db00d8;
mem[8] = 144'h00c60285036a00fc02100268fd3b001103bf;
mem[9] = 144'h00e201f3026003260352ff1bfe2ffde30347;
mem[10] = 144'hf74ffd21ff18fcdcfad0014efe8ffd9dfe8b;
mem[11] = 144'hfdb300dcfec9003001c800f6fd71fe5a0219;
mem[12] = 144'hfd73fa06fd9c02dc00a9fb10fea3ffd6fe4a;
mem[13] = 144'h010d027a009701e4007f026f02b901060023;
mem[14] = 144'h007a00dc03910363027aff93fdae01af02cb;
mem[15] = 144'h01f20435035702f500dafd85fd30feb3009f;
mem[16] = 144'hff40ff5c0159007600b4005dfec2ff040079;
mem[17] = 144'hfe5d003affa2fe460163ff67fee8ff6fff05;
mem[18] = 144'h0069ff62fdd8fdf301800036ffc0ff1a007e;
mem[19] = 144'hff90ff39005bfdec0113fff0ff8cfeaa0013;
mem[20] = 144'h0121006dff06000effe3fdf6ffb8fe170108;
mem[21] = 144'hff2f00b8ff3c005c0052ff1dfeaa0103ff42;
mem[22] = 144'hff71005fff4ffe6701dcfec8fe2c0119fee2;
mem[23] = 144'h00660096fe8900f2ffea00e8011e0073014c;
mem[24] = 144'h00e1004efedaff8cff580089ffca002400b3;
mem[25] = 144'h003bffd80079ff8b0082010bffc700db0057;
mem[26] = 144'hfec4ff81fe2fff4b01b1ff3eff450086ff2a;
mem[27] = 144'h015400fb00eefeb5007bff8600b60081fef3;
mem[28] = 144'hffb4fffffe1affda0037ff6eff5200f5ff7c;
mem[29] = 144'h017201590176fef600fcfeb5ff06fdc20001;
mem[30] = 144'hfe960099fea3ffb6ff04010401bc00ea0235;
mem[31] = 144'hfef4ff71ff000073fff8fea900effde300fc;
mem[32] = 144'hfebefecd016600c500a000bbfe07ff49ffe2;
mem[33] = 144'h0171009eff3b01ddfebdfeb8008dfe37ff3b;
mem[34] = 144'hfe5efe320073019fffb50058ff59fff9012b;
mem[35] = 144'h00f8005c00bc00540048ff96fe590025fe46;
mem[36] = 144'h00defe51fdfc00870152fed80134004f00f1;
mem[37] = 144'h00ad007300e0ffcf01d200cdff64015d01d1;
mem[38] = 144'h00bbfdd4fff8fe3801b1fec0fffb0032feca;
mem[39] = 144'h0029000c016b014100bafedcfedbfe5ffe23;
mem[40] = 144'h00cdff3a008aff69fe35fe64fe35ffcc0186;
mem[41] = 144'hfe0cfe1dfe4bff6afeb6ffe7fe250073fee2;
mem[42] = 144'h000dfe3e011bfe88ff31fe7b00a70184fe9f;
mem[43] = 144'hff06ff1300f300e4ffc4fe7d005d0161ff5a;
mem[44] = 144'hfec8ffa1ffdd00e3007cff3b00adfef1fff5;
mem[45] = 144'hfe3000d40105014f00d6ffc6ffea006f0160;
mem[46] = 144'h000a0153012b014ffe6f0071018bfe660157;
mem[47] = 144'hff0c0090017700ccff38018cfe11fe81fee2;
mem[48] = 144'hff02feecfeafffe1fd76000f01010080001b;
mem[49] = 144'hfe5fff5cfe7600a40056ffcd00fafdd9fffa;
mem[50] = 144'h0053ff48000dff55010aff2afdca00b4fe79;
mem[51] = 144'hfdf9feedfeefff17ff7fffe7ffd1fec6fd6e;
mem[52] = 144'hff86002cfe8afe11feb6fe6dfda6fd58ff35;
mem[53] = 144'h0094ffbdfeeefe31ff28018b013cff79fe97;
mem[54] = 144'hff0dfebc0045012600d70092ff6d000700bd;
mem[55] = 144'h0046ff0eff42fff0fd730074fdfb00f100f6;
mem[56] = 144'h010ffe8dfe5900fe0082fe0ffe1dfe94fe6c;
mem[57] = 144'hfe07fe8cffafffceff2ffea400d4fe0100af;
mem[58] = 144'hfd9bff1e000100670110fdf8ffd7fed5ff9a;
mem[59] = 144'hff00ff02ffb400d8fde3ff70fe15001aff64;
mem[60] = 144'hff2eff02ff74fff7fdb1fdaefe1affd9ff5f;
mem[61] = 144'hfe25fdeeff5b00bffe5500e1fdf800b6ff9f;
mem[62] = 144'hfe3fff90fddb0038ff1c0082ff2cfe13fffa;
mem[63] = 144'h004dffa4fdeffde5ff810068fe530082fd97;
mem[64] = 144'hff51fc00fec5fda6fdcdff02ff88003b0453;
mem[65] = 144'hfb0ffcc10341ff80fe5100a9ff7e046a009f;
mem[66] = 144'hfa81035cfd41018c009ffca1fc800219ffa3;
mem[67] = 144'hfe0ffe3701feffccff7001fc01880468ff63;
mem[68] = 144'hfc71fcf0fcebfb71fe0bfe3eff41016e035c;
mem[69] = 144'hff8cfd92fee201c50185ffedfff4fe6cfe81;
mem[70] = 144'hfbb2fbc6031bfef0fe0000ce009304c70320;
mem[71] = 144'hfec4fce0ff8affbcfe0600de0171014f0141;
mem[72] = 144'hfd05005201d4fe99fe61fd92ff0f019801ed;
mem[73] = 144'hfa6cfd99015bfe47fc9bfef9ff2004230324;
mem[74] = 144'h06f700ebfe93ffd500d2ffc2fdc4fb57fe39;
mem[75] = 144'h018afe28ff0c017c011000f2015bfe660142;
mem[76] = 144'h002707000330004a008002e3066004260099;
mem[77] = 144'h0293febafa89ffd9fe57fae2fd36fd31025e;
mem[78] = 144'hfc3ffc2c02dfff37fe51fed200fa00c9011e;
mem[79] = 144'hfc49fa3effc1fdf6ffcafea0ff7203b00318;
mem[80] = 144'hfdef0163003c0148fdd6011e0025ffaefe64;
mem[81] = 144'hff06fe5b015e01cbfe81fe4a013600f60026;
mem[82] = 144'hfffc008aff3aff23009bfe1b000000d70003;
mem[83] = 144'h009600370175fdc30159fe42fdf2feb801cc;
mem[84] = 144'h01750163fdbdfe310159ff00ff14010b0116;
mem[85] = 144'hffcb00d4010bffa8fef1ff91ff9bff15017c;
mem[86] = 144'hff73fe36fffc0020fe2d00cbfef201360096;
mem[87] = 144'hfe41febafe4e007f01a0ff0eff9900e900ff;
mem[88] = 144'h01ae017cffedfe03fedb0057fec3fe41fe59;
mem[89] = 144'hfe0fffe9ff44ff1b00370011ffee000100f5;
mem[90] = 144'h00c9ffc9008701260086fed0ff630121ff43;
mem[91] = 144'hff980221ff8d0070feca005900e8fe67feaf;
mem[92] = 144'h003c00b8fe16ffb40079feaefff30222fe05;
mem[93] = 144'h01f2fe0aff9ffee20169013900b3ffe4fe7a;
mem[94] = 144'h00acfea10105013a00a2ffd8fe8f01c6ffd1;
mem[95] = 144'hff66fdfdff93fdc1003a00c7ff64ff55018b;
mem[96] = 144'hffe603920514ff5fffa1047a045104ea046c;
mem[97] = 144'h0278064207cefb23faf1fdf3032bfe5eff75;
mem[98] = 144'h04bd06090179facaf7cbfc460082fdbeff68;
mem[99] = 144'hff3902040331000802b5fdaafe9e01fcfec7;
mem[100] = 144'h015701d303cd0060ff230134020f01e2026a;
mem[101] = 144'h007b008202e101e9019c01c3ff87021a0105;
mem[102] = 144'h005d03cd0a0cfeeefd47ff4a015903e9fe6e;
mem[103] = 144'hfff9027601cb01a9fec30274ffdb017f01e6;
mem[104] = 144'h0556076807f0f7a5f9c2ff5f02aa00b3fff9;
mem[105] = 144'h0231068e05edf883fab6fe4401980121009f;
mem[106] = 144'hfa7afd4ffd9c00f7fd79fa90fd6e019e022a;
mem[107] = 144'hffe7fdec031cfffffceafd09fdc0013901b1;
mem[108] = 144'hfe1c0197fde7fdeffe4bfba1f6adfd4afeba;
mem[109] = 144'hfcad0058040d024a0637065505ca056b0557;
mem[110] = 144'h02a106b4072dfd38fcdafd57fef901520079;
mem[111] = 144'h029603f00778ff1efe3efff5013f027e00dc;
mem[112] = 144'h00b0ff4e008cff1e01eb00ffff02fea200cf;
mem[113] = 144'h0083ff7d0161007d007a01a50076007a011b;
mem[114] = 144'hfe6300b4008500e3fdf801bdfed90137fdea;
mem[115] = 144'h00ac0088ff0d0155ffb60057ffabff68ff18;
mem[116] = 144'hffa50175fe8b00c4014afecb00ddfefdff50;
mem[117] = 144'h0052002c011bfe2c0161fe8affd0fefc0051;
mem[118] = 144'h017400030162fe040178fdd9fec000820114;
mem[119] = 144'h01a9010ffed6ffd40072015a007bfe2a017a;
mem[120] = 144'hfe7600a3ff0efefeffc8fee1ff71fe8efe79;
mem[121] = 144'hfddc0138ff1cfee10004fe19fef50163fea5;
mem[122] = 144'hff8aff08008e017f0005000efed1fe80fea3;
mem[123] = 144'hff65014f00f0ff07ff5dffc9ff63ffbc004b;
mem[124] = 144'h00c4fefc012efe16fe98fed8ff84fe47ff66;
mem[125] = 144'h015a002dfebffec2004bfe1400b10057ff72;
mem[126] = 144'hff370060ffcb01b200500109023affc00106;
mem[127] = 144'hfe56ffba010fff0cff150105fef700080023;
mem[128] = 144'h00c6fe88fdc5fb0efefe01a80097fe59fac4;
mem[129] = 144'hffcaf9dffb08016f01b401ce0254fcc5ffff;
mem[130] = 144'hfd9afb71fe180052fff9fbb10048023d0098;
mem[131] = 144'h006602edfd9c0034007d023702b40185ff83;
mem[132] = 144'hfccd00d0fda7fd220091ffcc01f2003cfd4a;
mem[133] = 144'hfe870002fe1e014f001e022900780040ff73;
mem[134] = 144'hfecaff0ffa25fc65feb0000d00d2ff56fc7a;
mem[135] = 144'hfeeefed5fe53ffeafea4006102540134fd6c;
mem[136] = 144'hfff1fc46fbae011e00f1ff7e00a4febffc32;
mem[137] = 144'hfdaaff3bfc0301ceffed02940470fef6fdb3;
mem[138] = 144'h028903ae02fa02d4ff3bfce602100284ff6e;
mem[139] = 144'hff4f01e2ffd500e5ffbefe3101be02a4fe0c;
mem[140] = 144'h03f704f603980016ff7a061b0218fe5901dd;
mem[141] = 144'hfd25fe80fff0fbeefb55fd58fd2ffcf7fb3a;
mem[142] = 144'h015dfd6df87fffa6febaff1a0313ff65fe50;
mem[143] = 144'hff5bfecdfe2afda5ff8400c00199005ffd70;
mem[144] = 144'hfe1101e9029403c1027901740027ff7402c1;
mem[145] = 144'h0298fed500a400aa0281059802e20085fe8c;
mem[146] = 144'h025dfedcfdd0ffde035b0ae506350198ff8d;
mem[147] = 144'h02bd01e4022700cf00b0ff71ff9fff43ff6a;
mem[148] = 144'hfe8dffb200ea038a01fa0344000f00d3fed6;
mem[149] = 144'hff57023a028a030803bdffa2029f0091018d;
mem[150] = 144'h00d40151020a040b00f70191023e00e9ff37;
mem[151] = 144'hfeae00640267042b0188fff301d6ff74ffea;
mem[152] = 144'hfeeb00a501d103a8061a04a003d7feda0135;
mem[153] = 144'h001a0190016703f104fe041c040bffea00a1;
mem[154] = 144'hfc0501af0088006d01b5ff69035dfecd0061;
mem[155] = 144'hfded02ab00d400fdff6e01620147001801d4;
mem[156] = 144'h04dd0153001eff8502dd029f01210139002c;
mem[157] = 144'h0012032f034f042600c2fe77fd0a0124014d;
mem[158] = 144'h02990311033f04e9041e007503cbffd60220;
mem[159] = 144'hff2a005602f8032001a1021e00e1feb700c7;
mem[160] = 144'h01bbff68ffe3fd45ff3efd91fb09fc250174;
mem[161] = 144'hff65fb2701b80057054c0146fe78035f03fa;
mem[162] = 144'hfa2c0251ff84042a064907260517034e01ab;
mem[163] = 144'h0225fae8035cfcc7fe21fe02000705bf01f8;
mem[164] = 144'hfd18ffbe002f0013ff2e00d4fbbdfe3c017b;
mem[165] = 144'h0306fe22fea60062ff4c0061fef0fe92fe5e;
mem[166] = 144'h00a5fa65ffc5fe5eff1101b9ff84ffb3038e;
mem[167] = 144'hfecfff7dfea2fe77ff4bff85fd9efc460071;
mem[168] = 144'hfcd7fc8801df02d703bc0287ffc9019f03c9;
mem[169] = 144'hfbc8faa301d1ffeb001efebefee8ff53024b;
mem[170] = 144'h00f9047affa203be00a408f80637ffe3ff12;
mem[171] = 144'h0149004afe6001b5fd680130ff3afe24ffea;
mem[172] = 144'h028b044b036eff69031701f405b8081c021b;
mem[173] = 144'h06840406ff54006bfe66ff50fed9fb09015a;
mem[174] = 144'hffebf9bc01d2fd84013c03b2fe38005d0231;
mem[175] = 144'hfe64fca701fafe07fee801bdfe2200390285;
mem[176] = 144'h0176fdddff500055017d00bd0158feb9fe51;
mem[177] = 144'h0104002eff5fffc3fe1effa2010e001901da;
mem[178] = 144'hff94ff73fe13ff20ff1401b6ff0bffc0ffb0;
mem[179] = 144'h013afea9ff81001efed5ff3b020000e0ff15;
mem[180] = 144'h000afe4afecdff24013101adff990176fef7;
mem[181] = 144'h01860058ffaffe88ff82fe3d0005014a0061;
mem[182] = 144'hfef400cbff0e00ac013bff30ffe7008cff3c;
mem[183] = 144'hffedff87fe8aff79fe7d0141fed7ff58fe69;
mem[184] = 144'hfffd0236fdf3feb1013500a2fe4afddafeef;
mem[185] = 144'h009fff9e011cff4dfef601320007ffda018b;
mem[186] = 144'h0094ff0b0178fe9f0041010efedbffa8ff4e;
mem[187] = 144'hff6bfee7ff31ffab0013000d0014ff6bfe15;
mem[188] = 144'hff61ffe600aefe5afeacff17fe62fff70100;
mem[189] = 144'hfe29fef9fe81009f0214011dfecd00f10036;
mem[190] = 144'h01920177001e01970043fdf0fe6dfe21ff84;
mem[191] = 144'h00ea00c50028fedd011ffe74fea3ff08ff47;
mem[192] = 144'h026effadfe48febdfeadffb101cb00f00058;
mem[193] = 144'hfcebfe22fe33fd7efc4afc87fe5afce0fc7f;
mem[194] = 144'hfb8f01b0ff560067f8b1f556fa02fca8fe07;
mem[195] = 144'h00a8fe70fec900d600e902e8028efc4bff60;
mem[196] = 144'h002b0025011cfcb600a4012b037700ad0063;
mem[197] = 144'hfe470103fe2dff75fec3feccfef7fffb00c2;
mem[198] = 144'hffe7fed6012f00abff8f002efff9ff0dfbed;
mem[199] = 144'h0079000800a8ff45fe67003d0112fe58fdcc;
mem[200] = 144'hffa20079ff58fe49fdb00015fe02fac2fbfe;
mem[201] = 144'hff4d01f2011dfd12013501fbff95fc48fcd1;
mem[202] = 144'hffc9fff300d200e1fdc6f9adfea0ff2bfdde;
mem[203] = 144'hff7002050072fe9c0208ffd00315ff87febf;
mem[204] = 144'hfc8efdadffe500d1fdb6014ffcddfce30064;
mem[205] = 144'h00d5ff2c0002fe56fe3afe8802910129ff71;
mem[206] = 144'hffc8fdf4001ffdc40013fee9fe4bfd21fc81;
mem[207] = 144'h013efecaffa2ffde01d50224022e0003fe86;
mem[208] = 144'hfebcfa59fa92ff72fec5fbf2fcd3fffdfd57;
mem[209] = 144'hfb60fcefff41082805d502befcdf0308018b;
mem[210] = 144'hfa1c037a004a0332086b046201dc02ed021a;
mem[211] = 144'h01cafd870386026efe1101df07da051d03a2;
mem[212] = 144'hfdbbff25fd97fff603d9fe96fc7800810297;
mem[213] = 144'h0002ff77feaffdef0134ff44ff16fdf7fed6;
mem[214] = 144'hfc26fae6fe1802370404ffef00f2fe8e038b;
mem[215] = 144'h0104ffb3fe25028a022cfdaf0088000c0215;
mem[216] = 144'hfcb7fd50fbd408c30680ff62ff810115008f;
mem[217] = 144'hfb83f9a9fbd4065e03fd0001ff71023004a5;
mem[218] = 144'h09f7036b0077026d06300b0000bbff06ffeb;
mem[219] = 144'h05330069fce2024e05fb05e902100115005a;
mem[220] = 144'h06d006890114064c02f103fb0ea2051e0168;
mem[221] = 144'h03e5fe90fd2cfd53f990f6f1fb79fbfbfe9a;
mem[222] = 144'hfc61f8fdfe3303770545023800c9023b032c;
mem[223] = 144'hfd5dfb94fcb804070386fee0ffbc02d802a3;
mem[224] = 144'h0079fea601c203b300f60158ff260132043f;
mem[225] = 144'h016300d504d8ffe700ab08fe032f01b40255;
mem[226] = 144'hfe9202ee008100f502d0066d0055019700ec;
mem[227] = 144'h031bfec300e3031800d10080fe8f032c0060;
mem[228] = 144'hfc9f012200c4fe0c01020411031afefa0310;
mem[229] = 144'h01ab0061ff9001d0ff86ff4b0122ff8b0141;
mem[230] = 144'hff6b010104890062ff1102e903d5037501b4;
mem[231] = 144'hffbbfd00ff66ffa4ffc100ac021a0192019a;
mem[232] = 144'hfe27ffff02fafcaa05af0a6204de02c00263;
mem[233] = 144'hfea1000e024afc92023107ea067a03600435;
mem[234] = 144'hfd07fe68fe1c018bfe6cfde501fbfd59ff9c;
mem[235] = 144'hfd23ffb3fdfffea8ff450154017dfd6802a5;
mem[236] = 144'h0181ff72028300a3030c01dcfd4003780026;
mem[237] = 144'hfddf0015fc35039c0086fd89fd32fee200e2;
mem[238] = 144'h003effc00550009a00ff059b0316030dff9a;
mem[239] = 144'hfe00ff7f02b1004dfef6046f0203013affa1;
mem[240] = 144'h02970362ff190004007d0382032affb4ffcb;
mem[241] = 144'h054dfe55fa4b01e7019bfef4008800e20262;
mem[242] = 144'h0156fbb7ffae031e024bfd9d01f802bd048f;
mem[243] = 144'h034f034c02adfde1001f02f3ff08ffd10003;
mem[244] = 144'h0092012bff4e0395fd90034b0247029d01b2;
mem[245] = 144'hffc0007501d1ff5301ac00de013b00e10084;
mem[246] = 144'h059c00bdffae0059014f00360187000000d6;
mem[247] = 144'h043c019701a00231feb9017200bb00fb0087;
mem[248] = 144'h02c8fd0f0026ff70ff91fee2ff2200b7009c;
mem[249] = 144'h0266018bfe91fdf2ff18ff5d0197010cfeeb;
mem[250] = 144'hff82033e03c4013efca7ff6b01bd00f903bc;
mem[251] = 144'hffc2009700420307fced00ed01ca0248fff3;
mem[252] = 144'h026105610346fd7c028b010bfd4401dd029e;
mem[253] = 144'hfda7fe1c003b017701ab0317046b0018017c;
mem[254] = 144'h055f00b0fc91fd500154ffb5feaffffcff21;
mem[255] = 144'h04a20265fd53001dff0401a501f20103023d;
mem[256] = 144'h045a03b4008701c00136027b02f50300fcbe;
mem[257] = 144'h056801fef974fec1fe4b04e7033dff110023;
mem[258] = 144'hff7bf79202770036fe500345ffe902cd037f;
mem[259] = 144'h02dd0757fcafffd3fee90259ff55ff41fd05;
mem[260] = 144'h01ba065102fd0089016f0138027d0089fe8e;
mem[261] = 144'hff9a014a0057fffcfefcfcdc00630097032f;
mem[262] = 144'h04d304d2fcc2ff6f010d0146015b023efdb6;
mem[263] = 144'h015c0287030b02cd002402ed0183ff27fe4c;
mem[264] = 144'h03a20168fdb8fdd1fe14058c02b4fdf6fdda;
mem[265] = 144'h02b602c9ff4ffedafe2105190285ff5ffe7c;
mem[266] = 144'hf62b01b5014301a1fb42f6f300c2048c0087;
mem[267] = 144'hfeb905ee05680070fde1fa3d019701fe006c;
mem[268] = 144'h0251005f0107ff1efddffe37f624feee01c8;
mem[269] = 144'hfd15002bffed0292053d041d050703830094;
mem[270] = 144'h04ae02b8fb57ffb50002015d0327fe6cfd09;
mem[271] = 144'h022e061c00d30099ff10038c03c9fec3fc67;
mem[272] = 144'h03c002800261fe76ff9f012901de02640562;
mem[273] = 144'h03e904f70414fd10f9b0fdf1fdc3035800ec;
mem[274] = 144'h019302630448fd5ffbb5fda0009d01800293;
mem[275] = 144'hfff90175fe20fedd02ac0092fb860150ff22;
mem[276] = 144'h02c800bd012f0124feb3002cfef2ff7e02a3;
mem[277] = 144'h042a014a00830174021d0147021b014f0239;
mem[278] = 144'h01f5032c03b3fcbefeccffd4fd19022c003c;
mem[279] = 144'h02a0000a033affe5fe9a013dfe57ff020379;
mem[280] = 144'h0323027e046bf961fadd006200e2026d01cf;
mem[281] = 144'h024103470304fae4fa2fff40ff2dff1000e5;
mem[282] = 144'hfbd7fd6dff7c033bff53ffbbff4dff3f0303;
mem[283] = 144'h0054fdef026eff6bfb58fee0fcfffc9403c3;
mem[284] = 144'hfbf7ffaf00bbfbfbfdc1f9c6f78d01020183;
mem[285] = 144'hff5a03430312022b03f006d5040600d4050e;
mem[286] = 144'h02060360056cfe49fe82fdc5ff3a009800c8;
mem[287] = 144'h03e1034a02affe39fd1affb5fea7feca001e;
mem[288] = 144'hff48ff7500d0ff6a027600d300ef00b20210;
mem[289] = 144'hfe7afd35ff5d009e025e0434065c0295fe20;
mem[290] = 144'hfd45f9ee0089fdfa00ea07e0012dffa80274;
mem[291] = 144'h013e02c8ff8d0145004101e004dc0702ffec;
mem[292] = 144'hfe79021d028701fb000a021b024300590337;
mem[293] = 144'h0019fef600b901d7fff6fec3fdf9fff20254;
mem[294] = 144'hfe63ffc60042010e01ba037002bb06a2ff67;
mem[295] = 144'hfee5ffed003b001200f3014f001003370258;
mem[296] = 144'h005802ffff6ffdfa0439058b01c0fff70131;
mem[297] = 144'h00a4017e038500710136041202b602dc0121;
mem[298] = 144'h012600ea0063ff3dfe7afd96fe8c01cc01a9;
mem[299] = 144'hfd74010100b900e4fdbefedf00a6016a0267;
mem[300] = 144'h05490782046c01a4ffe9007303c702dc00ec;
mem[301] = 144'hfd51fd4cfc8901840328fc7dfeba01acff8e;
mem[302] = 144'h0141fe21fe21fe0f006d02b102ac05a2fe44;
mem[303] = 144'h010001ea0149fe59010d043d03b301c702c5;
mem[304] = 144'h0042ff900099ffa500be00d4fff8fecfffd4;
mem[305] = 144'hfdca0134fe94fe2afe8ffdd5fefe0156ff5d;
mem[306] = 144'hfe5dff9200c6ff07ff180133fe31ff13005d;
mem[307] = 144'hfe4a017100e8fe1ffee80063ff4900f9ff51;
mem[308] = 144'h01450056fe46ff98fe7300ebfe9afeadff29;
mem[309] = 144'h01cdfed301d90026feec0043fe7e00adffa0;
mem[310] = 144'hfe72009d000aff10fef9002c0155ffbdfe2c;
mem[311] = 144'h000000bc0044fe4efe43fe4cfe8700fdfe02;
mem[312] = 144'h0009feabfffaff1e00a8ffdcff370036002e;
mem[313] = 144'hff5dfe0d0076ffabff2aff9900e2ff9b015b;
mem[314] = 144'hfec9fe86004bff7e007eff1cfe3400230045;
mem[315] = 144'hfe60fdaeffa0ff98ff65006efdccffc4fded;
mem[316] = 144'h0133fe2eff300039ff79fddc0109ffd000cc;
mem[317] = 144'hfd790116ffa1ffebffab0069fe490063fe80;
mem[318] = 144'hfedc018d010100e7fde7ff8cff0aff26ffc8;
mem[319] = 144'hfdf700800091fe7dfe6efe0900e00130ff2c;
mem[320] = 144'hffdffdeafb1d0150ffc300dffe05fcbefc5e;
mem[321] = 144'h01eafda8fc13062805b8ff45fcdffdaa03ed;
mem[322] = 144'hfbdcffec0285048a090e0196ffc3021a027b;
mem[323] = 144'h02c7ff98fdb1fed7028c03c504ffffd302cf;
mem[324] = 144'h0051fffafd4b0332ff4efe09fd3afee1ff37;
mem[325] = 144'h001bfcb1008f000ffedeffeffc520069fe27;
mem[326] = 144'h00b4fed1f97900110310fff2ff79faab01c8;
mem[327] = 144'h0015fff7fd3601eb01bfffa3003d0070fdf1;
mem[328] = 144'h015efb6efa5f07de033efa05fc0eff4f0089;
mem[329] = 144'h0019fcb1fae904f802a1fc85fce400b7febc;
mem[330] = 144'h03f703100299024e0156053601500207ffba;
mem[331] = 144'h02be0129ff7701fb04d601f6ffe90203000c;
mem[332] = 144'h01c6ff2001c3017103cd0166067402bf00ee;
mem[333] = 144'h009900f3ff4dfcbcfc23ff710234ff6bfc76;
mem[334] = 144'h0082fe97f98a03e1042fffcefed9fbf80062;
mem[335] = 144'h037c00e9fc6e02020080fee4fe7efee60055;
mem[336] = 144'h01feff2bfeb5fadafb4dfea90336fd41fde1;
mem[337] = 144'hfd8afc83fc16fe80008bffe0000bfc2dfed6;
mem[338] = 144'hfc8cfbc700ef0093fd64f98cfd9a02880104;
mem[339] = 144'h017400ecfee5fdd3fdae053a0317ff160032;
mem[340] = 144'hfec1006d0085ff5ffcebfffc025202cefd00;
mem[341] = 144'hff21007e000a00c4006d019b00bd00d100c1;
mem[342] = 144'hff88ff00fa89fac4ffca024a0144fe8afcdb;
mem[343] = 144'h02ec03260050fed6ff96ffd702fb0020fec6;
mem[344] = 144'h01aefe84fc5efecefe69fd33ffa5fedafc23;
mem[345] = 144'h010a0112fbb0fe2ffeb7ff1b03f1fde4fc8b;
mem[346] = 144'h04db041d01e9025fffd5fd670204011500e8;
mem[347] = 144'h00440314007e0187018fff8f042601470119;
mem[348] = 144'h034d0320fff100fbff4505090179fd0502ad;
mem[349] = 144'h017fff6dffe8fcdefc19fdab021901a5fdf8;
mem[350] = 144'h00acfc3efb13fef6fe2400bb0045fecefcdd;
mem[351] = 144'h0058ffd7fd48ffb1fd850046039affe3fd67;
mem[352] = 144'h0134004b0452002cfea5fd35ff1cff980078;
mem[353] = 144'hfe04007701cffefefc3df9c9ff0aff16fe2a;
mem[354] = 144'hfdcd023fff90ff97fe7a032f02b2ffdd00e5;
mem[355] = 144'h0276facb02a40047fe4dfa7302c7fe9f019b;
mem[356] = 144'hfe3c023d012afe9bfd85fe7bfc64fea6ff52;
mem[357] = 144'h0113ffcdfd5eff6d004201d2002cfe7dffa6;
mem[358] = 144'hfe3cfd3501c700cefd04fcffff39fc73004e;
mem[359] = 144'hff3700ab0172ffe2ff9bff5efc79007aff65;
mem[360] = 144'hfe87021801f0fc69fc1df896ff34fd35fda3;
mem[361] = 144'hfcaeff0f007afe7ffcacf92efa51fdafff8d;
mem[362] = 144'h031e0164015f008e0602073aff5300d500af;
mem[363] = 144'h00b4ffd200aefefd039a04c3fc60ffe6fea7;
mem[364] = 144'h02adff0100b901ecff73fccb0447013e01b5;
mem[365] = 144'h047c031302fc035b052601f1ff3a01470273;
mem[366] = 144'hfe2afe0802a0fe2dfdc0f9dbfdb9fc460259;
mem[367] = 144'hfdddfe53023f0193fd79fd63fc7dfde7fe76;
mem[368] = 144'h00ea01540004010bffd2ff63018dfe2300ee;
mem[369] = 144'h0192018d01b4ffaffe57ff70ffd400a20099;
mem[370] = 144'hff81002dffc501ad0069ffb000abfffdffd1;
mem[371] = 144'h0050ff1a0034008effc0ffcd006bff6dfe95;
mem[372] = 144'hff3dffffff69ff50fe780038ff1efeabfe86;
mem[373] = 144'h01a8fe750038019ffe5a01d001b900bbff3c;
mem[374] = 144'hfe03ffdf0072ff61ff9600bb008cfead0039;
mem[375] = 144'hff7a00e5ffa300b9ff3fff10fe7eff4a0196;
mem[376] = 144'hff67012800fe0134fe80fe59ffe90021fe8c;
mem[377] = 144'h0042fe1e003400e8fe86ff3e0185fe21fefa;
mem[378] = 144'h00f70000014cfe660042ffb3ff4900050073;
mem[379] = 144'h01220158fe88fec3013600ae011100970003;
mem[380] = 144'h001f00dcffc4fe02ffe0fef1fe990009014d;
mem[381] = 144'hfe00ffb0ff31006bfff101b0017300240115;
mem[382] = 144'hfeb700bafe97ff29ff79005aff9a01bdfe8d;
mem[383] = 144'h00f60167016ffff9fe7efe07ff03ff55fe25;
mem[384] = 144'hfeb9ffbcfe6afe63fee4fd61fd4600f500ae;
mem[385] = 144'hfef5fef5fddffe2cfedffdddff140123ffdd;
mem[386] = 144'hffbbfe6100b30000fe8c026c01edfde6ff6f;
mem[387] = 144'hfe27fecafdf6fe82fff5fe21010102770245;
mem[388] = 144'hfe3afe48fd6100e7fdf1ff40fe02013800fa;
mem[389] = 144'h0122ffb2fff9feb100e2fe510002feec0025;
mem[390] = 144'hff00006dff9effa8fdbfff67010800660309;
mem[391] = 144'h0004007300a9ffbbff82ff6efdb5fe3801d6;
mem[392] = 144'hff0bfda3ff3300890003fea50067009400b5;
mem[393] = 144'hff03ffce0097fe7dfe990038fe2fff7b01cd;
mem[394] = 144'hffeefedcfe9b010501b100b3fd21ffad00b2;
mem[395] = 144'hfd6b004c0113fde1fe22fee6fcf900e6fe5f;
mem[396] = 144'hff47026700c1fe90fe21ffeafece006cfdce;
mem[397] = 144'hfd53000c0091fdd7febefff2fe90ff10fdeb;
mem[398] = 144'hfe92001efd78ff66ff86fd8bff8300ce0255;
mem[399] = 144'hfd85fe57fdcbfeeafd83fdf1004fff18ff6f;
mem[400] = 144'hff06fd900219fdf0fd4efa55fbe5fd5f00bd;
mem[401] = 144'hf978faea037f010f0150fe16fd89004b025a;
mem[402] = 144'hf742025200c8010e095d074704420240fe5b;
mem[403] = 144'h0214fa1b0367ff1dfd3efcb0023004ab01fc;
mem[404] = 144'hfd58fdabfe7fffd8ff6ffd33fa8efd0a0095;
mem[405] = 144'h0261ff78ffd6febe02900177ff1bfe11009f;
mem[406] = 144'hfcaef86e017bffb2fca3febefd5800aa0286;
mem[407] = 144'hfd2cfea7feb50184fd83fbe6fd51004d0182;
mem[408] = 144'hfacdfc28ff3d03c30425fd2afa20ff0902d0;
mem[409] = 144'hfbdefd18003f00ebff48fbf6fc2600cb0144;
mem[410] = 144'h06e40450fd80028008ba0c3900bc0007fd5c;
mem[411] = 144'h00c7fe30feed012903d10438fe5affbdffc1;
mem[412] = 144'h052b0269043a00a9023a03b10c6404c60309;
mem[413] = 144'h05e901c7029bfcdefc6cfbc7fb0afddc007d;
mem[414] = 144'hfd4bf8f7022101be0029fd41ffbffe310183;
mem[415] = 144'hfe40fa56ffaffea1fe09fb17fb27002c0385;
mem[416] = 144'hfb7dfcafffbbfe97fd75010dffcaffabfebd;
mem[417] = 144'hff89fe49fc6601b700bf00780055ff9dfce6;
mem[418] = 144'h0129008afec5fe40ff0800daff5bfcf1fc85;
mem[419] = 144'h005fff16fe19fe8f001d009afd6bfd96ffde;
mem[420] = 144'hfcd1ff49fe1f00d0ffdb018dffe3ff46fce3;
mem[421] = 144'h00eb017efe5ffe21ffa5ff450072ff0c018b;
mem[422] = 144'hfdf8fe30fe4cfc5f01670109018efdbaff97;
mem[423] = 144'hfe6bfe99fcdeff9afd200075ff77ff12fdb6;
mem[424] = 144'hffcafdfbfc39013affdf01f7020e0068fdeb;
mem[425] = 144'hffaefe82fe55011cfe42008902030049fd25;
mem[426] = 144'hfcf5004ffe51ff4afbb8ff34fe0dff84fddf;
mem[427] = 144'hfd9bffb8ffa0ff35fbe6fd36fe3b00ac0032;
mem[428] = 144'h0255ffdcfd44fec7fe32ff1ffc7bfca4fec8;
mem[429] = 144'hfdc2fb7dfc0cfe39fddbff4dffa5fcf1fd54;
mem[430] = 144'hfee5fe26feceff78ffd200a20336ff11ff54;
mem[431] = 144'hfeabfdf4fe6c0107fdbaffc80026fe49fcf6;
mem[432] = 144'h01420048fe37ff9ffe82fffafef9ff99ffd6;
mem[433] = 144'hfe200115fe8f005bfe540031001dff55fe28;
mem[434] = 144'hfffdfe7a003cfe3cfe3d008d0090ffa8ff8f;
mem[435] = 144'h007d00ac0134fe3fffe6fe820130ff8cfe8f;
mem[436] = 144'hfef3fdee0099ffd6ff6efed90159ffbd0139;
mem[437] = 144'hfe8e0156ff5d00d8006efff7ff9bfecaff47;
mem[438] = 144'hffc5fdd1ff6cfeb3ff17ff230143ff5e00ce;
mem[439] = 144'h0071021b0059ff79ffc2014dffd701c0ff13;
mem[440] = 144'hfe2fff19feaaff81fee4ff9ffdf4ff64ff7f;
mem[441] = 144'h007cfdecfdcb01ef00cefeabff4900680033;
mem[442] = 144'h0086fe6afef6008dffe0012aff9e0027fe60;
mem[443] = 144'hfdbefe0000640091fe7ffe0f0064fea9ff03;
mem[444] = 144'h009301650160fe8e0148fe6bff26fe44fece;
mem[445] = 144'hfe93fdfaff6e00d400fa00e600a00053ff40;
mem[446] = 144'h016d010c00bdfeda0121ff2a0110006f0000;
mem[447] = 144'h00e9ffb5fdcbfee800baff33fe82fdde00b4;
mem[448] = 144'h00460030ffbafeba0077ff20fefffeb7ff41;
mem[449] = 144'h001000140010ff1a01d10168016dfeef01a2;
mem[450] = 144'hff29fe2dfdeafec2fed9013500d8fe6f00bf;
mem[451] = 144'hfdbdfdde0047fe6cfe4bfe1effb5013efeee;
mem[452] = 144'hfeb5fede0143014f00cd00df0096ffb5ffe4;
mem[453] = 144'hfea500e4ff9dff3cfec9ff8500d6000901e0;
mem[454] = 144'h0070ff79fec1fe64fe570105004afe81ff61;
mem[455] = 144'hff41ff190066ff0afe35000afecaff31fe8e;
mem[456] = 144'hfeaefe0100670060fe67ff9f0024fe170138;
mem[457] = 144'h0170006cfed2fe9a020bfee8fe650088ff68;
mem[458] = 144'hffd1fe9dfea8fe1bffcdffacffbafe40ff75;
mem[459] = 144'hfecfffa8ff5c0063fe2c003ffed60014ff70;
mem[460] = 144'h0090fe6bfe1d008afeb0ff16ff9bffb100e3;
mem[461] = 144'hfece00b4fe9d001c00b5feb30175fedffe8a;
mem[462] = 144'hff93ffe600e7febf010b0182ff370139ff12;
mem[463] = 144'hffb8fe74ff5f016e0146fe71ffd6fff70179;
mem[464] = 144'h0397feea0321fef70059ff46010afd340123;
mem[465] = 144'hfbddff4203abfd21feccfc2bfbe00036fd38;
mem[466] = 144'hfed60253fe53ff37facef9b6fe1bff2ffe1a;
mem[467] = 144'hfcc3f955ff5bfeb70092fff2fb8dfdb300c4;
mem[468] = 144'h02d3001f0030ff6cff11fe49007efce0fd4d;
mem[469] = 144'h000a01050046ffe9ff800118ff0e00920146;
mem[470] = 144'hff5dfd7d01bbfdd401a90004fcb6fd90ff8b;
mem[471] = 144'h031c00630085ff68fe66ffddffedfcb5001b;
mem[472] = 144'hff82febb03a7fc7bff7800ccffdcfe21ffb2;
mem[473] = 144'hfedfff96ff81fe53fe7200c40165feb4fde6;
mem[474] = 144'h0184fe13feca001400f4fe4d01de000efe54;
mem[475] = 144'h0247ff99fe2aff6cff25fdb30198fef6fd52;
mem[476] = 144'hf85af741fde9ff01ffa50119f6ccfb45fd7d;
mem[477] = 144'h0281020400abfe8ffed500000230fe93fff6;
mem[478] = 144'hfba0ff230428fea2ffd200aaffb7ffe501bc;
mem[479] = 144'h00e5fece0174ffa2007d001afe29fe3dff19;
mem[480] = 144'hff3dfcbb03b1fe5eff20ff26002d033b03d9;
mem[481] = 144'hfbe204bd03fb015bfcf5fd2e01b900d900df;
mem[482] = 144'h05820750ff810014f910fa480081fbecffdc;
mem[483] = 144'hf99bfe35010500e303dc001e00ae020d00f4;
mem[484] = 144'h0286fdc8fee2fed70175ffc7020301e200cb;
mem[485] = 144'hfe84fdcafe37fea8ffa50242fef6fff3ff75;
mem[486] = 144'hfd39001a0246ff640227fec8fe8b01eb0092;
mem[487] = 144'h0153ff5dfe9301a800ea028d0116024affcc;
mem[488] = 144'hfe930530028dffa4fbdffefd0541fdf700c0;
mem[489] = 144'hfe4800e201ccfef1fdc100750257036500d6;
mem[490] = 144'h018effeafe36000e009f0034fe8f0147ff93;
mem[491] = 144'h02fefc79fd1e02c805650390ffbc03ac0175;
mem[492] = 144'hfec70026ff62002b020501c2fd63fcc300c2;
mem[493] = 144'hfd96fbd101e9fd5c005d0024033801890120;
mem[494] = 144'hfb78ff15037a01d10029ffab010602230121;
mem[495] = 144'hfefcfe87023c00f3ffd8ffe3ff6a01550278;
mem[496] = 144'hffd3ff4a00000148fef1008d001d001500fb;
mem[497] = 144'h004c011b0093ff49fe77fef3fe600161fe3d;
mem[498] = 144'hfeb7ff21ff5b0104fe68fe20000400d80088;
mem[499] = 144'h011f00e4ff3ffea900a20095ffacffb9ffc4;
mem[500] = 144'hfef3fdf4ff85fddeff37fdb90105ffe1fdd2;
mem[501] = 144'hfe5d0037015901cffe39ff00ff5fffdb0136;
mem[502] = 144'hffde01fefff5ff60004fffcbffd3fdc20191;
mem[503] = 144'h007f0159ff3f019bfeca00dffe6bff8cfff5;
mem[504] = 144'hfe53ff18ffe2ff1d0127ff80fefefef7ffb0;
mem[505] = 144'hff8ffea70022fec900b6fe5b00f4ff7bff20;
mem[506] = 144'hfe62ff8a006f0042003a008e000600ad00ac;
mem[507] = 144'hfddcff80003fffe6feedfe4eff34006700ee;
mem[508] = 144'hfdd300d9ff33fe2e008dffb60092ff23feba;
mem[509] = 144'hffcafe03fea10067fe3fff80ff6c007c013e;
mem[510] = 144'hfed2ff18ff08fe450064fe6c0091fe3ffdd1;
mem[511] = 144'hfe25ffbc00a4fde800cc0007fec1014cfe69;
mem[512] = 144'h004efd6efe4bf8b2fc1dffc201fd012bffb8;
mem[513] = 144'hfe3a01e70392fdf9faebfc6703f0045e017a;
mem[514] = 144'h01af023002080259fed6fe4bfeaffdddfe2d;
mem[515] = 144'hfe0ffe1eff0ffa7efed001eeffdafffe0154;
mem[516] = 144'h0028ffabff39fd65fc72fd80fffb035b0121;
mem[517] = 144'h0205fec600ba00a80009005b002affc1fea6;
mem[518] = 144'hfcf3fd7a0267fbf5fcdeff9d01df025f039c;
mem[519] = 144'hfef1fe7c002efc35fe1ffc6b011d0159009d;
mem[520] = 144'hfdb20329fe67fe0bf93aff180477021e00c8;
mem[521] = 144'hfd0a012a0134fc13f9e0fbab018704590296;
mem[522] = 144'h0447ff60fdd600f804400293fd0d016cff04;
mem[523] = 144'h01ff0052ffac0339ff0300c601600435ffbf;
mem[524] = 144'hfe6aff8dffa3fdffff1804230317fe5ffede;
mem[525] = 144'h0337fe9201c6fc88fca9fcd4fdf301a000ce;
mem[526] = 144'hfb45ffb60148fe14fe62fc3001e00597037a;
mem[527] = 144'hff2bff82fff0fb36fbe9feaaffa50184007c;
mem[528] = 144'hff62fd220120fff901d0003d00de0089034d;
mem[529] = 144'hfedd00da00ba006f02e7043d066e05c8ff64;
mem[530] = 144'h0128fe55fe9e029002f50871056a035400a7;
mem[531] = 144'hff9a039805b90135fe6a013302ba08f00229;
mem[532] = 144'hfbe400ad0108fe77ff8101b203a20190016c;
mem[533] = 144'h011e00b80186019cfe600043004101eb021d;
mem[534] = 144'hff70ffb5ff320071ff1a023c04aa05b40108;
mem[535] = 144'hfe36fe7500d500510168ff4d0225030f0229;
mem[536] = 144'hfe6e00ecff8e004301ad064905f9067a02ab;
mem[537] = 144'hfbabfe89ffe9fec50006030f034f0436054d;
mem[538] = 144'h04a4014d015802af0264fec3fe84fece019e;
mem[539] = 144'hff0801dc01d7ff10006cfffa038402af006b;
mem[540] = 144'h02300a9e0529015b02940496034a048e0074;
mem[541] = 144'hffccfb77fdb30131ff9afc01fa90ff32ffe7;
mem[542] = 144'hffd8fe5a006dff00002d045004df065eff0c;
mem[543] = 144'hfc4afe0f00d0002e02910104041b05f001f0;
mem[544] = 144'hfdad013bfeecff37fdcc013800a10024007e;
mem[545] = 144'h004cfee4fdb3ffe2ff77ff60ffdbfeab0019;
mem[546] = 144'hfea2ff1bff14ff7bfffe006bfeedff78ff26;
mem[547] = 144'h0150fe8e0125fffd00f8fe96fe50fe8d000a;
mem[548] = 144'h00bb003efe17fdf8fe3bffde00eeff5900b3;
mem[549] = 144'h0057ffa1ff68fecbfe460142ff65ff390016;
mem[550] = 144'h001c011fffcdfe79febdff5bfda8fe70fee7;
mem[551] = 144'hfe75ff67013affd7fe9fff150097fdadfe42;
mem[552] = 144'h0061ffbafeb9ff81fff00016013bfe3dff5e;
mem[553] = 144'h0148012aff15008cfe800022ff50ffa0ff50;
mem[554] = 144'hffc8fe3cfda3ff87fee2fe6bfdadffc2feb4;
mem[555] = 144'h00d9012f014600e200d80138fe1cffc2ff41;
mem[556] = 144'h0078feaeff29fe05fecdff1afe14ff3c0003;
mem[557] = 144'hfe04ffae0140fdc5ff18ff7c0130fe9a0092;
mem[558] = 144'h00d7ff0bff8efdf6fe4efd9e0074fdfcfeb8;
mem[559] = 144'hff700047001cfe41fe7001490037ff7cffe2;
mem[560] = 144'h006603faff1d060604b002340077febcfe1b;
mem[561] = 144'h03760072fafe0235045d069e038802e5fe10;
mem[562] = 144'hfe6af7f90062007303b30912021601bd003c;
mem[563] = 144'h04f50608ff6f01790107005ffdbe0284fe0b;
mem[564] = 144'hfd1200c5016f01e702630112003bff000075;
mem[565] = 144'h0190ff0a0162ffb90279fd5603000025ffb1;
mem[566] = 144'h014d0271fe5101af0313050503020392fdbf;
mem[567] = 144'hfd590089ff9a01a101510210017f01adff1c;
mem[568] = 144'h0293fce9fec703700684074f02a702f5014d;
mem[569] = 144'h01f60087fe77027604cf05710463fffdfeeb;
mem[570] = 144'hf84d029eff78ffa4fba9fb5a012801260014;
mem[571] = 144'hf94002740367fe4e00c301ae0323feec0059;
mem[572] = 144'h01d600fe00bdfeca0020ff8eff8302a7014b;
mem[573] = 144'hfe88004efd6903500296fc8bfd19fdc0fe8c;
mem[574] = 144'h013e010cfce801e4028602d2035302a4fcb0;
mem[575] = 144'hffb2012eff7b023b0445039a03570032fe4d;
mem[576] = 144'h0148025f018b010e009a043f0359fde60052;
mem[577] = 144'hfeabff93fc85fec5034103cf01afffaaff04;
mem[578] = 144'hfda2fcfbff15febcfd1cfea3fc7c02d8ff1d;
mem[579] = 144'h027001dffe5e028f01cf00a3fd73fd7dff48;
mem[580] = 144'hfabd0163002dff360216020c020cfda0fef5;
mem[581] = 144'hff06fe27009d0033ffe400f8fef00110ff06;
mem[582] = 144'h02fcfee7ffef01b100f1026f02b8ff4afd43;
mem[583] = 144'hfd63020000bb00f3fe7c02550068fe65ff30;
mem[584] = 144'h011300abff51009e022a08490085ffc30134;
mem[585] = 144'h0104fed500e2ff2e04110407023aff02ffaa;
mem[586] = 144'hfc460079feefff2afbc6f812ff72fd3dffba;
mem[587] = 144'hfdc5015a0146fdd0ff50ffcd0418004aff11;
mem[588] = 144'h014afcb0fe59ff4101c4021cfb88ff4cffb9;
mem[589] = 144'hfea302230110ff0e002ffb4efe61fdd20093;
mem[590] = 144'h0026fe04fc2201a200fa020403a7fec2fe36;
mem[591] = 144'hffd600f8ff12019401ac04a7019dff17fcea;
mem[592] = 144'hfe59fe28fe76009cffc6feb2fea9fe34014b;
mem[593] = 144'hff2c00f201cb012c01980033ff5f00cffe3d;
mem[594] = 144'hff750102fe7601d6fe88008f01010157fdaf;
mem[595] = 144'h00f5ff3b015d00c5ff96ff7cfdecff2aff6f;
mem[596] = 144'hfef000f9ff88ff9001b90046ff590114014f;
mem[597] = 144'h00ae00e0ffb0ffe6ff14ff3a005801a10172;
mem[598] = 144'h001f00abfe66013d0102fed30074002aff8a;
mem[599] = 144'hff5101d90064016ffe84fea0fe7afeb60190;
mem[600] = 144'h015fffc80114fe0fff83fdf9003afe89ff75;
mem[601] = 144'hff63ffb5012b016e022afde80072fdec0031;
mem[602] = 144'hfeedfe7f012afe1d00faffda0036fe22ff18;
mem[603] = 144'hff10fdcd0117fe4cfe36fdbd001cff4bfe40;
mem[604] = 144'h014bff7f002aff1300f800e80018ff74ff42;
mem[605] = 144'hfff2fe25fe11febaffd80138ff4cfe68fdc8;
mem[606] = 144'hff72ff71ff2600020079ff20ff0d00da00be;
mem[607] = 144'hfeb500bbff8afdd5ffffff9efdfdffbeffed;
mem[608] = 144'hff08ff4900d60226ffc600df010f01180286;
mem[609] = 144'h022e0073027a011103c7050404e2061e00eb;
mem[610] = 144'h039f028800200279062a0d330a8703d5021e;
mem[611] = 144'h03a0fe8e02cffec4fea3fdc90189010b060c;
mem[612] = 144'h018bffd5ffb804ef010afd89fee7010cfff5;
mem[613] = 144'hff880191fef90115ff43fef4fe8c01ab001b;
mem[614] = 144'hff46ff4102a1004fffdb00e802f501bf0475;
mem[615] = 144'hff9c010effbb039c0083fdb2ff3600a700a8;
mem[616] = 144'hffcffee7029d02d103b304cb02470360ff81;
mem[617] = 144'hff78004b0046028201de033100ca027a0006;
mem[618] = 144'h0194005801b50265032102eefec200670166;
mem[619] = 144'hff4202820017fe6bfcc6fd64ff39008e0224;
mem[620] = 144'h01f90300028dff12fff1ff7c01df019a0072;
mem[621] = 144'h0490fedefee7ff1402a4ff3f0055003b025f;
mem[622] = 144'h0088000000c2ff33027401bf045e04250272;
mem[623] = 144'hfeb5ff09ff9001db0101fecb00260147018f;
mem[624] = 144'hffcdfe7f0156fff4fedafe2afea90071ff12;
mem[625] = 144'hff9100acfe55ff46010d01affebd003aff1d;
mem[626] = 144'h000c023dff22ffb900c40066ff860178ffde;
mem[627] = 144'h00370013ffbbfe05ff2efede01ecffc300bf;
mem[628] = 144'h0061012bff34014500a1fe130061fe71fed8;
mem[629] = 144'hff5dffe8fe6900e7010f01acff6201e1003c;
mem[630] = 144'h0081007afe1afed0020a0103022d01ceff4f;
mem[631] = 144'h00befe98006cff55ff12fe0bff42ff0f0167;
mem[632] = 144'h013effd5ff6e0046febf0015004eff80017b;
mem[633] = 144'hffeb004600d20097fe5eff71010a0048014f;
mem[634] = 144'h00910088fedf00f2ff0fff9401a001460040;
mem[635] = 144'hff580138fe5fff0a0112fede00d5febe0029;
mem[636] = 144'h0120ff06013eff69017cfeadfe22019ffecb;
mem[637] = 144'h00000009ff84fe6b014cff1a014ffead00d3;
mem[638] = 144'hfe9b015a017e00d4fe9e01bd00a500f600e8;
mem[639] = 144'hfdc8008000a00135010dffb800c700990116;
mem[640] = 144'hffaa024a0514063704a9006b01bc003c01d5;
mem[641] = 144'h02db035501de0266022102c102f8fc82fef2;
mem[642] = 144'h038702f2fda5fdeb0019084b016efadefec7;
mem[643] = 144'hfd8fff4fffc106800221fcd70098feafff03;
mem[644] = 144'hff0e0123026302c1037b02850106018fff2c;
mem[645] = 144'hfd31ffddff1affe9fe92fecb01dd0201002d;
mem[646] = 144'hff290126041d0604008f005701d8ff380117;
mem[647] = 144'hfe91ffff03c6057d04c6fff80234004cfe1e;
mem[648] = 144'h002303a80232014902a203a000b5fbe3000e;
mem[649] = 144'h013301c603fa024d042a02e70053fe81fe82;
mem[650] = 144'hfdc8fe2dfe5cfe80015301de001efed6fe4e;
mem[651] = 144'hff1cfd9b02befe97032101b8ff59ff37fdf2;
mem[652] = 144'h0076fd24fcb10051fdeafef1fd61fcd1006a;
mem[653] = 144'h01a50332057504400651014600a2027b0253;
mem[654] = 144'hfed802ca027c0479ff7400a60131fd8a0102;
mem[655] = 144'h00f200e50507057c028b01af032700aafe9e;
mem[656] = 144'hfe9200940061fe8afebb0189fe24feb7fe04;
mem[657] = 144'h019701bd0054018800bc01ccffa000f9ff52;
mem[658] = 144'hfe65015b0152020a0166ff50011bffe0ff9a;
mem[659] = 144'h01e0fe6800a7fe710010ff8effdc001bff1c;
mem[660] = 144'h016e0082012b0033ff6efdb9fe44fef500d9;
mem[661] = 144'h0038ffca0174fe71ffa2fec6010cffdeff83;
mem[662] = 144'h00e7024cff05ff26016b002e00a1fe3cfe8c;
mem[663] = 144'h00ef012900f30067ff98ffce0051fee3fea8;
mem[664] = 144'hfeb5fec2011c001afe93fec90099006cffae;
mem[665] = 144'h003dfda60144007a014e00aefee4fe2500bf;
mem[666] = 144'hff4c00aa012efebefe90feaf001bfe4d00ec;
mem[667] = 144'hfdc7ff0ffef2003300bbfdd2fec300b00178;
mem[668] = 144'h00fc00dd0022ff9affa900c8ffeaff94ffdd;
mem[669] = 144'hff56fdfffe05fe20ffeb015700f3006efe8f;
mem[670] = 144'hfee9ff89011efea4fe70ff37fe86fe0d007a;
mem[671] = 144'h00b8ff97fe3eff0bfffffeb2fea8ff19fecc;
mem[672] = 144'h02390254fed003870132ff03ff85fd08fb6f;
mem[673] = 144'h00adfa83fb360504053a04a50230ffc70289;
mem[674] = 144'hfca3fc98fea103a4076408b405bb036f0078;
mem[675] = 144'h060cffbbfdbaffe9fe3400480250fe2ffed2;
mem[676] = 144'hfd620145ff76026801f1ff3ffec5ffa0fee8;
mem[677] = 144'hff7e01b301b900e400e8fe4000a0ff59fe67;
mem[678] = 144'h04570062fab502f9010c04610137fc8bfe5f;
mem[679] = 144'hff1b00ec00f301ec02dfff25feafff50ff2b;
mem[680] = 144'hfe64fdf2fb6106b7078901340072ff3cff63;
mem[681] = 144'h00eeff64fb8405a206bd035a01aafd70ffe1;
mem[682] = 144'h015002f303cefe5c02800604030800f30054;
mem[683] = 144'h0018025f024bffb2ffee0377032effe2fd08;
mem[684] = 144'h03a400020031006c02f604b8035204a3023d;
mem[685] = 144'h031304e00137ff4ffed1fe5ffd4ffd13fe7c;
mem[686] = 144'h02bafe66fb400275030e03d0014bfdfffec9;
mem[687] = 144'h0116fd84fcda00bf040b03c50140fd65ff29;
mem[688] = 144'h03ca006e032d02f4001afeb4fbaa02980287;
mem[689] = 144'h0108034a07b903ac00c4000b000e01670100;
mem[690] = 144'h02060984007bff240727065101aafd5afe9e;
mem[691] = 144'hfdd7fe8d02650399ff3afdb0fde003960345;
mem[692] = 144'h033c033500ee022801c5fc47fdde0121010a;
mem[693] = 144'hfcd9006cffe4ff73ffdefce6fbec005fffd8;
mem[694] = 144'h0020013103e2031b010fffccfef8005d0433;
mem[695] = 144'h023a0145ffdf023201e5fdfffc63008300bb;
mem[696] = 144'h02520222050404ad045cfed0006002a905fc;
mem[697] = 144'h0177017401cc01570102fe92fd0b000d03db;
mem[698] = 144'hffacfe31fd54ff49023a059702b100890164;
mem[699] = 144'h03f8ff73008b01550326ffdefd89ffbe0276;
mem[700] = 144'hfc56fc9800a702590172ff630496042dfea6;
mem[701] = 144'h04730050002e00b2017efe54021f019e0347;
mem[702] = 144'hfd7701b005e001f502530153004403be05d0;
mem[703] = 144'hfec90266024c009fff89ff1afde6ff4803f6;
mem[704] = 144'h0434033901cb000cfda30081fed203a20691;
mem[705] = 144'hfd7c03280572fea4fdc4ffdbfeb2fec9fedf;
mem[706] = 144'hfa61035c02d3ffe0ff9b017bfb0dfd20fd2f;
mem[707] = 144'h002bfd05ff41fde6ffbbfd23fcb104f2febb;
mem[708] = 144'hff7203880291ffb7fffefd5efea1fdd803ee;
mem[709] = 144'hff2bfd9afe59ff6dffa0fabdfd99fdfd0025;
mem[710] = 144'hffe500f70301fe0efea001a6ff260382001d;
mem[711] = 144'h00fb030e03dafdbffce4ff38ffbdffbb024e;
mem[712] = 144'hfed903fb0394fd0c015901dffcf9009503ba;
mem[713] = 144'hfe15043f0602ffe2ff3f0099fc59fe9902cd;
mem[714] = 144'hfa8afdfbfffe0023fd24fef2fd97fccb0013;
mem[715] = 144'hfd8f02750305fecfff02fe46feebfcd4040c;
mem[716] = 144'hfae2fc09fb61000efe13fc70fe0d0200fda9;
mem[717] = 144'h03c1004d0008ff0bfd8400f8003303d00448;
mem[718] = 144'hfec501ab0681ff8bfd48ffc6fef001bfff3c;
mem[719] = 144'h0003032103e6ff8bfdfe00ccfe68ff1402a2;
mem[720] = 144'hfdbafdf102adfed50298fe9fff6901f404a0;
mem[721] = 144'hfda90160040e00cbfbc70063069406be0150;
mem[722] = 144'h03a50213001cfebbfe6c00ce05ffffacff62;
mem[723] = 144'hfdd40216054501620031ffd001f6047e013f;
mem[724] = 144'hfd80ffed0112fe5b024501f604460542005b;
mem[725] = 144'h014a02a800bb026ffe69013f0426ffd5fe73;
mem[726] = 144'hfce4ff630450ff99fde9fe0a0344056302d3;
mem[727] = 144'hff07ff1a021502be001b0000022504170072;
mem[728] = 144'hffe10030fffafe83fbfa0182060c021e0096;
mem[729] = 144'hfedb00d50263fe34fd89022704c606480130;
mem[730] = 144'h04f101f2fe0101f0050e012afd9fff620125;
mem[731] = 144'h0334ff70fde30298047c02f401d100e30273;
mem[732] = 144'h013306410312001dfd5d03410539fff7010e;
mem[733] = 144'hff2dfab3fd7a0082028dfc9dfe48ff2e003d;
mem[734] = 144'hfdb0006103710107ff2c00c403250716007e;
mem[735] = 144'hff30fe790376ff76fec8012e058a04e203fc;
mem[736] = 144'h00f9009ffeb200b400540176feb5fe7d00bc;
mem[737] = 144'h0067febf009e00ba01aeff00ff0900eb0033;
mem[738] = 144'h0133fdf60010fed4fe35fe52ffb9ffa800b7;
mem[739] = 144'hfff8fdc70074ffd5004801410028feb10183;
mem[740] = 144'hffe3009b003cff23ff9c0012fe3cfee8fe6f;
mem[741] = 144'hfec901dffe7afec6004500e4ffd4fe83fecb;
mem[742] = 144'hff9500610080fdcdff0d0107ffde0175fed4;
mem[743] = 144'hfedbff8b0075009500ff00e6ff400064ff26;
mem[744] = 144'h015cfed1009eff15010a0147ff7ffe490077;
mem[745] = 144'hfe4b0178003700a9fec401b601c80028fe75;
mem[746] = 144'h00cafe4e015afe69017ffe6600800082fddd;
mem[747] = 144'hfec90033ff2a003cfe86008dff92fdf40012;
mem[748] = 144'hffcbfeeafde6fe10feb6fdec0120ff0d00de;
mem[749] = 144'hff60016f012cffd100af017bfee8ffe3ff68;
mem[750] = 144'hff2c01c8ff9201a7fffcff6affbc0169ffa8;
mem[751] = 144'hfeb9fe2900af004100d7fe4d00e4000b0117;
mem[752] = 144'h01210049016f0557fff7017203ee006bfe06;
mem[753] = 144'h005a02d50045fdb3fc7cff0f0066fbb2fe3c;
mem[754] = 144'h026b014ffe7afca8f9fd0037fdc0fd1afea9;
mem[755] = 144'hfcbdff4affcc052cfef602ca006dfedc0014;
mem[756] = 144'h0023ffa702f0ff60ff1aff2303e1029afe0f;
mem[757] = 144'h00fe01430121febd00a000eeffdb0170022a;
mem[758] = 144'hfec2020d0128012ffd4cffd5004afbfafff5;
mem[759] = 144'hff0f011e015f0394004200e203c7019ffdf9;
mem[760] = 144'h00f2029d00defe0bfc70ffdf0321fc01fce0;
mem[761] = 144'h0291022d01b400d4fe8c00600344fdb9ff30;
mem[762] = 144'h02f0fee000e800da0468007cfde10381009d;
mem[763] = 144'h00bcffc8ff16ff250558005b0174036cfeb8;
mem[764] = 144'hfc58fd3efd790111fe8d00d5fc75fd0201a0;
mem[765] = 144'h010f00b30459071203a9011f00330310ff27;
mem[766] = 144'hfda4ffc903eb0136fb97ffa4014ffc210111;
mem[767] = 144'h0005004501be0206002702100278ffba006a;
mem[768] = 144'hfedcfec5026102b80172ffe1fdf0ff19024f;
mem[769] = 144'h011701840718fff9fdfcfed9fc79ff1402ae;
mem[770] = 144'h03ad07a400440160fde8fd14ffc7000f0061;
mem[771] = 144'hfec9fae7007b02d901e8fee7fd55fb81024f;
mem[772] = 144'h02ecfe98fe6bfff401c6004700d500b400e7;
mem[773] = 144'hfea2000cff3e00d2ff780158019afe2afeff;
mem[774] = 144'hfd79ff48026effbb02dc014000c8fc3c01fc;
mem[775] = 144'h00ccfe7e00db009100d5ffabfffdfefefe44;
mem[776] = 144'hfe5b01f00320010300a0fe2a02e2fc54fe38;
mem[777] = 144'hfe6dfd25ffd600dcfe3ffc39fed4fe7effd0;
mem[778] = 144'h026bff78ff51ff60030705ce00c0feeefe4a;
mem[779] = 144'h04e4ff1fff15ff860309026e0027fe130013;
mem[780] = 144'h0032fb89ffed031a019a025d00d1fc05ff7a;
mem[781] = 144'h01ca050a06fa000900d80347022001d10267;
mem[782] = 144'h0023009a040b016a0189fcf6ff05fc730388;
mem[783] = 144'h020afef10138ff5d01e5fdb3fe74fef00110;
mem[784] = 144'h03a402e201320137fe87012e025804520619;
mem[785] = 144'h0101058807d8fe28ff24003601b401ddff5c;
mem[786] = 144'h0020048c023bfd2e02780779fe13fef500f1;
mem[787] = 144'h0114fe7cfef600effedbfffe01760541ffec;
mem[788] = 144'h028704e603e8fefb00fbfecafe5302c103b8;
mem[789] = 144'hfd04fee1fe66ff46ff66fc2cfe2bfebf00c4;
mem[790] = 144'h016c035103ebffc4fedeff74004104af016d;
mem[791] = 144'h00e60113041c025000af008d003e00ea047f;
mem[792] = 144'h026e085503b1fd70008603a3fe3c045d0524;
mem[793] = 144'h0425052c065800450045ff46ff43025c0633;
mem[794] = 144'hfe9b002f002b024c003d0110003902d80041;
mem[795] = 144'hffbf00d201cffed8fe39ff94ff78ffed04ed;
mem[796] = 144'hfcfbfe2100a80122ff97000cfee3012bff59;
mem[797] = 144'h032fff74feb8027d017f01430426062a0509;
mem[798] = 144'hfeee02400423008aff1202b8ff1303d4017a;
mem[799] = 144'h01de0311042001170018ff3afe59046703c7;
mem[800] = 144'h005cfe5000c1fdadff37ff8a0040fdbbfff4;
mem[801] = 144'hfdfdfe07fee8ffdfff6dff00ffb5ff16fd8c;
mem[802] = 144'h005fff65ff01fe0ffe9a009bfdc9001dfd61;
mem[803] = 144'h0016fe53009a004e002d00520060fd77fe66;
mem[804] = 144'h003aff5bff7dfe4efd9e00a60093000bfdb9;
mem[805] = 144'hff37011600f9ff2a00bf0012ff4e00e1feed;
mem[806] = 144'hfdeffe01014aff90fda0fedf008eff6700aa;
mem[807] = 144'hfe8ffedf008efe66ff65009efdcafe41ff6e;
mem[808] = 144'h005ffe9afd53fe12fe5e00340079feb50101;
mem[809] = 144'hfe40015ffe20ff0f0028fe68fe6e007fff1b;
mem[810] = 144'hff58ff05feef0058fef4ff34fe370191fdd1;
mem[811] = 144'hff31fe7efe86005ffdeaff590078fe930094;
mem[812] = 144'hfdfdfff5fdb2fdbf007cff39ff68fdfefe91;
mem[813] = 144'hfe2b014dfee7ff16fdc2ffc9ff6c003ffe72;
mem[814] = 144'hff36fe24006a00a7ff31fdddffad017cfdf9;
mem[815] = 144'hfef5fff90055ffe1fdeafe95fe75fdc601a6;
mem[816] = 144'h02600306fc15017a021cff7cff4ffad3fa9e;
mem[817] = 144'h02e5fbd4fb0a0393068a00ecfea2feb302c2;
mem[818] = 144'h00abfda9fe8901d508fc07ef0416022c0178;
mem[819] = 144'h03080071fea100f0ff630105ffabfe310234;
mem[820] = 144'h03f60174002702470406fef5fee1fc1afd37;
mem[821] = 144'h01540228018f005a0118fe15013cfe63ff6b;
mem[822] = 144'h0201ff7ef8d7040003770087008ffbe300cb;
mem[823] = 144'h02c10280ff4e0182034901cc00feff44fc7b;
mem[824] = 144'hff49fde3fa4b092805f4ffac008f008d000c;
mem[825] = 144'h0323fd72fb8006ba0517ff3ffeb1fe2cfe60;
mem[826] = 144'h033801e1030f00880057059303fe04640199;
mem[827] = 144'h03ff01b902d2000304b3ff28035401ceff44;
mem[828] = 144'h03a8ffb3ffbe0509016aff7e036c01d303f0;
mem[829] = 144'h00d9063f01700193fdd101cf03eefdf7fd1c;
mem[830] = 144'h0312ffecfaba04120284008bffdbfea90132;
mem[831] = 144'h03e9ff8cfd890369038d0091fe36fd94fed4;
mem[832] = 144'hfe63fe1afcf8fa95fe8c02990155fba7fe4b;
mem[833] = 144'hfddbf9d5fbd2006afee5fd5cff40026a0358;
mem[834] = 144'h0135fdd5fe8003f1ffe5f7b6fddc04fafffe;
mem[835] = 144'hfc0f030a024dff8cffd00238012e00db026d;
mem[836] = 144'h0108feb1fcebfdcf00a500c2002400a7fd80;
mem[837] = 144'h007100fafe4f011d0134fe4fff0bff8d0179;
mem[838] = 144'hfda6fc78fc73fe1fffe301b4012fffa3ffd9;
mem[839] = 144'h00d1ff4efdfffd0100d6025c0224ff740042;
mem[840] = 144'hffadfd15fd7a017cfdcdfea100c7012b0034;
mem[841] = 144'hfdc8fc28fb49fffafe68004e0098017cfea7;
mem[842] = 144'h03bc03ad009d0171ff43fbe40197003fff6b;
mem[843] = 144'h0260002afe3302a30158001e01d800390036;
mem[844] = 144'hff4a0480030e02c8022905a700aa04c702aa;
mem[845] = 144'hfbfbfd40fdf3fac9fd4aff44008ffc0dfd8f;
mem[846] = 144'h012dfc31fbc6ff85ff9501f60051ffd0fed8;
mem[847] = 144'h0038fd91fbfafeafff2d009e008700d8ffc5;
mem[848] = 144'h01260334ffeefe4a0179024c0256fe12fd7e;
mem[849] = 144'h03c6ff8bfe430147004dfdf0feb401ba029e;
mem[850] = 144'h028dfd43ff5200c3fd4ffd0404b80513026b;
mem[851] = 144'h01f0ffee00a1ff0800e8ff62ffa6fc3b0123;
mem[852] = 144'h02f6000201b2fed2ffc0017001bffe4afe32;
mem[853] = 144'h0530028f001e0089007003c102bb011301ba;
mem[854] = 144'h031700c4008afd2d027300a00182000ffcb6;
mem[855] = 144'h00cc00cffffc0085002aff2500d6fe2aff0b;
mem[856] = 144'h01c5ff300154ff79003fff7e046501befe19;
mem[857] = 144'h04300138fe88fced0002003f009f009dfd6a;
mem[858] = 144'hffc2ff5b0251ff9dff3a0124028f03af0257;
mem[859] = 144'h01fa015801c401d1fc80fdfaffdc023700d7;
mem[860] = 144'hff5aff8802d10116fef50162fdd2fd8202d1;
mem[861] = 144'hfdc4046b028ffee701520381029a00270115;
mem[862] = 144'h044f005afddaffe8007400a8ffeefcc900c3;
mem[863] = 144'h0399022d0097fcd2000a00d9000afea5fe39;
mem[864] = 144'hff61009202c7016602b7053001c100bd03f1;
mem[865] = 144'h068403d604e6fca2fead00000208fd730157;
mem[866] = 144'h06d4052f009a0006fbd4fd610280015001ae;
mem[867] = 144'h02a4ff0bfe8302d4017b00e2ffb0fbec0077;
mem[868] = 144'h011c0188035901b3008d02df0089ffd0008b;
mem[869] = 144'h0220015e02ca018b0303002403ba03b001b1;
mem[870] = 144'h03140330038501e70142fe9fffbbfea4ffdd;
mem[871] = 144'hffeb01da0219ffdf02c102f200060181ffc9;
mem[872] = 144'h025202670347fecffca7001f02d901810213;
mem[873] = 144'h0226036104f3fed9fd27fe4e0222fd0cff08;
mem[874] = 144'hf9d6ffbafed9012d014e023c00890071028a;
mem[875] = 144'hff5dffc10058fe1dff86033fff40006c006e;
mem[876] = 144'h01c0fbcafd80ff8f029dff5ff8d4fb60ffcb;
mem[877] = 144'hfcfb01920254036d03e6041b03a2059a04ab;
mem[878] = 144'h02cf01e1067c014a01ddfddeff8cfe2600fe;
mem[879] = 144'h02370331024dffc200af01b502a4ff6bfe91;
mem[880] = 144'h0377025f0129041203db02e903c002710289;
mem[881] = 144'h03b6045a0433fc4b0027fdf8fc32febc0028;
mem[882] = 144'h007e05d50379fc89fda0fd84f9edfce3ff86;
mem[883] = 144'h008bfe4dfbf70210034c0009fe12ff33ff59;
mem[884] = 144'h011b02a50125ffbc00170280fe6f00c70508;
mem[885] = 144'hfec8ff8600770112007bfdff00f8fe300107;
mem[886] = 144'h03af022e01ff045b01ba01d2fd5c0122005e;
mem[887] = 144'h01c000af027a035f003dff81fef2ff700040;
mem[888] = 144'h05a6047d0568fd7cfd54ffa80099008003a5;
mem[889] = 144'h034a062a03590036ff94ffe9fe7701cb03dc;
mem[890] = 144'hf91afe05ffbdfef9fe920179ffd7fde5024b;
mem[891] = 144'hfdf6fe07feafff6bff5a01e0feb9017d046d;
mem[892] = 144'hfe4cf99afb23ffa0fecbfb74faf9fed7fd43;
mem[893] = 144'hff66034300bf05cd05ca04cc053a054401c2;
mem[894] = 144'h0345030303b00267ff40fee3fd2f02610211;
mem[895] = 144'h044c0178042e0338fedefffcfe4dff61ffde;
mem[896] = 144'hfd4efaecf7ccfaafffde0180fcd9f91ffb4d;
mem[897] = 144'hfecef9c3fcfa023401ce0213046007750323;
mem[898] = 144'hff8dfe2402c2031b018b031b073708130335;
mem[899] = 144'h01dafe210140fe1c005eff83fe32ff450395;
mem[900] = 144'hfccaff10f7d8fdeaff30ff5eff4afcadfe48;
mem[901] = 144'h0361000601ac0296018d03c504a301510307;
mem[902] = 144'h003ff956f8ccfd57019501f60248ffdbff2c;
mem[903] = 144'hff80fc19fb24ff39fd3b019100d8fe67fd0a;
mem[904] = 144'hfb82f927fabf01ad020204c402db036bffc4;
mem[905] = 144'hfe86f9d4f8c80038016903c00319021d0001;
mem[906] = 144'h073b04a600a8047c01a903160330025cfd6e;
mem[907] = 144'h01ea0091faae02be00df012604650034fc6b;
mem[908] = 144'h01a0030006e40359030801d2043c05d90570;
mem[909] = 144'h00abfde6fab4fcd4feeffd2ffc58faa8fa11;
mem[910] = 144'hfe87fbabf7d4fdb101b70068033c03ebff9f;
mem[911] = 144'hfe82f961f8acfe9f009f0300ffb4015c004a;
mem[912] = 144'hfe70fdf5ff0bff78fdb8fd76ff63fda4ffc0;
mem[913] = 144'hfebffefafe54fe6dff3ffea8fe76fee1fe19;
mem[914] = 144'h004cfe18fd9700f1fe9d00f8ff3ffd760066;
mem[915] = 144'hff3fff25007cfdc3ff4dfe44feefff89feb7;
mem[916] = 144'hff4fff4bff8d00090090fdcdfe5bfeaffebe;
mem[917] = 144'h001eff1dffbaff2e0196fe6b00d00004ff1d;
mem[918] = 144'hfeaafdca007900fcfdd0ffc9008100b500a6;
mem[919] = 144'hff04ff9bfe8a00b500bafe11fe5bfe47fddc;
mem[920] = 144'h007bfff1feddfe39002300adfe4aff32012a;
mem[921] = 144'hfde3fd90ff9efdfbff79fdb400e5ff7dfe8f;
mem[922] = 144'hfe6efe2e00bffd9afed4012701270068ffca;
mem[923] = 144'h000dfed8fe9400d5fefafebefe14fe4affc7;
mem[924] = 144'h005d00910017febefeb7fd930108fe41ffa4;
mem[925] = 144'h007bff7b004dff95ff24ff0cffd8fdfeffc8;
mem[926] = 144'h004f00d7fda7ff4fffec007afd96fe75ff00;
mem[927] = 144'hfe0dfe80ffcefed8ff12feff0089fe71ff32;
mem[928] = 144'hfdecff78fcd3fceffd820288028aff27ff4e;
mem[929] = 144'hfa80fe4cfdd8ff28fc9dff4a0061fddffe41;
mem[930] = 144'hfe0dfda8ffebfe7df887f2f7fc3dff70fefb;
mem[931] = 144'hff41fd5f0025fd13ff820298ffe90069fdb4;
mem[932] = 144'hfc870128fdeefe3ffe6300750161feff0077;
mem[933] = 144'h00deff8c0118ff47fe2dff82017c009cfed4;
mem[934] = 144'hfe5afb6300d5fc97ffcd024601140037000f;
mem[935] = 144'hfddd0058004efcaafcfc009e00dffe72011d;
mem[936] = 144'hfe9cfe910081fba9fd7a015d01e0fffffda2;
mem[937] = 144'hfe8ffdec0059fc6ffe410428032c017c000e;
mem[938] = 144'h020d01ea003100d6fccbf4880044fd8cfdb8;
mem[939] = 144'hff0800a7fe95008bfd47fdb60263fd9a00ce;
mem[940] = 144'hfe9e01acff41fe1affa9031bfc0201cdfdbb;
mem[941] = 144'hfd95fe2dff29ff05fbcbfc20fe08fd37ffa3;
mem[942] = 144'hfd80fd73fe64fc76ff1600e60284ff70ffe6;
mem[943] = 144'hfd64fcd000e1fda3fd8102450262fe86011d;
mem[944] = 144'hfdacfea3fe4bffbb0104009dfe52fd9d012e;
mem[945] = 144'h0029ff1c01590039fdf0fed5fef50042ff50;
mem[946] = 144'h00fa000d002000e5fd66ffbafe78ffeb0039;
mem[947] = 144'hfe6300760063ffc8ff150068ff3ffebcfeed;
mem[948] = 144'h003bff91fe11ff7ffdcdfe51ff7700350090;
mem[949] = 144'h00c0013201dbff63ffa3010000b700e7014b;
mem[950] = 144'hff3100da00730117006b0085002bfda1fe7d;
mem[951] = 144'h00d9fe14fdb8ff01ff17ffd20033ff67fe29;
mem[952] = 144'h0018fdf7019b006e00ecff59ff9bfdf5fdaa;
mem[953] = 144'hfe52ff4dff0cfd91ff97fe85ffa90013fdce;
mem[954] = 144'hfed2fffa006dfe7a006effc80039006ffdcc;
mem[955] = 144'h002efe10ffee0006ffaa0017fd9cff8f004f;
mem[956] = 144'hfffffe00fe3ffe08007ffff7ff3aff85ff4b;
mem[957] = 144'hfee2fe6afef20120fdf8004500b50037feb0;
mem[958] = 144'h00fd011001660022ff1eff1cfef50078fe9c;
mem[959] = 144'hfdeafdf2004e0131fe6dfe63ff1cfefe010f;
mem[960] = 144'hffc4fe990186ffdf00ce0165fe1d00ebfeee;
mem[961] = 144'hfe22fffbffbcfe49ffbdff4d00b2fe4a010e;
mem[962] = 144'hff15fefafe31fec600b2011ffdc6ffd3012f;
mem[963] = 144'hff38003aff5fff8300e3ffc9fe08fed80124;
mem[964] = 144'hfe4f0078ffcc000ffe38009efec80153ff1d;
mem[965] = 144'hff9bffec00c30032fee4ff30001dfee600d6;
mem[966] = 144'h0117feae00f3010cfe5ffdcdffadfe65fe79;
mem[967] = 144'h00620173ff5800f3011cffe501b901c8ffd8;
mem[968] = 144'hfea7009000f6feb1feec0146ff08006e0182;
mem[969] = 144'hff00fe5401080142fe48ff2afffe00c100e5;
mem[970] = 144'hfe2d00410162ffe7fdf5ff33014100dbffba;
mem[971] = 144'hfefafee7004dfdddffc6011000c8ff80fe1a;
mem[972] = 144'hfe6dff1ffef400c7ffa1fe3cfe4cfe0affa0;
mem[973] = 144'h00f1002100a50047002e001500b3fe8900b6;
mem[974] = 144'h012801d8ff7a00a101adfefb00dffec500a6;
mem[975] = 144'hfe47fea0019bfe16fe54fe32fec2fe53017e;
mem[976] = 144'hfd66fcc7fe77fe97fd4cffd8fd79fe19fdd9;
mem[977] = 144'hff9dfd31fe05fd13fdc70057003aff40fe35;
mem[978] = 144'hfef2ff57fe3cff2efe7000f8fe4bfe55fdde;
mem[979] = 144'hfe670241ff6cfe94fd6efef702be014000d1;
mem[980] = 144'hfd87fd29ffc9ffa9fdb7fdcd0044fd21fd46;
mem[981] = 144'h00200163015eff55010f0045fe230037ff7f;
mem[982] = 144'hfd2cff90fed0fdf9fed1ff760038ff6bff22;
mem[983] = 144'hfe50006ffd05ffcdfdbcfca10047fdb8012c;
mem[984] = 144'hfd4fff73fd3dfe13ff80fe720280003d015b;
mem[985] = 144'h005dff15fed5fd0dfce6fe30fffafee90001;
mem[986] = 144'hffed00150005ffe000a6fd04fe17fed2003f;
mem[987] = 144'h0095fdebffb7ffc5010cfeadfed8fe8a0079;
mem[988] = 144'h0126fdbeff1c0013ff41006501f3ff8e0071;
mem[989] = 144'hfe3ffe4dfe86fdfaff48fe5afe37feb1fcde;
mem[990] = 144'h0040fd94ff02fe5cfee6fdc90314ff370066;
mem[991] = 144'hff82fde30057fd1afd8aff310055ff9dfe27;
mem[992] = 144'h02ba02bd040603090108ff610016044b0374;
mem[993] = 144'h01f2068a053001bafe7dfde4fd47ff17fe81;
mem[994] = 144'hfd900736001ffed102a601e5fbcffa35fe5b;
mem[995] = 144'h0139fc12fe86ff7efeb7fe1703610145ff02;
mem[996] = 144'h043c045b01c401aa01a1fdf8fe1800d302c9;
mem[997] = 144'h0065002ffedfff90ff6ffc3ffda1fed1fe8e;
mem[998] = 144'h003701cd036bffb800effe8cfdf0fdfa0128;
mem[999] = 144'h01b4017102e2029e00e7fe2fff44ffcf033c;
mem[1000] = 144'h02450529057802c5fea6fda3fb6b00910473;
mem[1001] = 144'h036b054004e6fffe01b0fc4afc8d002c03e9;
mem[1002] = 144'hfe37fe4d018000d3028e04f4ffca01eeffac;
mem[1003] = 144'h03f8ff480218ffb901bf019dfc0bff130374;
mem[1004] = 144'hff62f917fc88ffc80011fe75007ffbfbfe9e;
mem[1005] = 144'h0390032104610202032d044c067d039d01d8;
mem[1006] = 144'hfecc02d804b9020a0213fe32fc7c004b0316;
mem[1007] = 144'h02ea029703be0326ff1ffe65fe84000a0069;
mem[1008] = 144'hfe63ffce01d00222010300eefe7dffeb0326;
mem[1009] = 144'h0121fcffff890493056a0376ff5e08250188;
mem[1010] = 144'hff7b013102b5031608300842077a044b001c;
mem[1011] = 144'h0269fe66022f01d90163ffb9fec605ce0355;
mem[1012] = 144'h009eff4d01b901c2010700c1fffefd140205;
mem[1013] = 144'hffbeff6a001b0090ffe1007a0210fe52ff4c;
mem[1014] = 144'h0210fe8b00e802ca012503d7fedd0347026f;
mem[1015] = 144'h0196fd5a005900c0026aff6cfdb50004035b;
mem[1016] = 144'hfe97fe140337059e05860494ff14037c0539;
mem[1017] = 144'hfea7fdee00c50425028d01c2ff31022504cc;
mem[1018] = 144'h03c601f2fff2018501aa097e0514007bffe7;
mem[1019] = 144'h003b02260029ffcefe0b034e01daffba0242;
mem[1020] = 144'h025c054601af0460011d0236060107ee0234;
mem[1021] = 144'h046d044afed80258ff17fed8fc0dfdfeff0e;
mem[1022] = 144'h025dff45012e014b01a5043b007f05d6045e;
mem[1023] = 144'hfe570052027f020d037c010efeb20042039d;
end

always @ (posedge clk) begin
	q_a <= mem[addr_a];
end

always @ (posedge clk) begin
	q_b <= mem[addr_b];
end

endmodule