`timescale 1ns/1ns

module wt_fc1_mem4 #(parameter ADDR_WIDTH = 11, DATA_WIDTH = 144, DEPTH = 1024) (
input wire clk,
input wire [ADDR_WIDTH-1:0] addr_a, 
input wire [ADDR_WIDTH-1:0] addr_b, 
output reg [DATA_WIDTH-1:0] q_a,
output reg [DATA_WIDTH-1:0] q_b
);

reg [DATA_WIDTH-1:0] mem [0:DEPTH-1];

initial begin
mem[0] = 144'h022e019d011d0453fea4fd2a008ffe86ffa3;
mem[1] = 144'h0083fefdfeb1fff0fd43faca0140fec60121;
mem[2] = 144'hfebcfc04fcad01100150fc0800b50423fd1d;
mem[3] = 144'h0150009f00180325ff73fcb400a5fff801b1;
mem[4] = 144'hfee9fe7d0039033501ceff0c0106fde4fd82;
mem[5] = 144'h0171010efee2ff8601c50194fe04ffd60000;
mem[6] = 144'h0072fec400c20189003efc4affe7feccfd57;
mem[7] = 144'h005d0027fc5402d6ff2bfff504b00278fc77;
mem[8] = 144'h00c7ff100135023cff6af9a902010064fef1;
mem[9] = 144'hfee9fe55ff9102de0287fcce00300041fc73;
mem[10] = 144'hfe75fc21fa05026800b200b1ff1dfa58efab;
mem[11] = 144'hfea4fc63fa3f03d900d00265fd2dfd72f7ea;
mem[12] = 144'hfdbd00f7ff870072f8a2fdbaffeffb05fdf4;
mem[13] = 144'h0066051208c3fac4fac1020a01a507b4062d;
mem[14] = 144'hff3cfed9005c0326ffaffab7032cffa0fe80;
mem[15] = 144'h00bdff7d005f03540230fdda00d70043fdc4;
mem[16] = 144'hfe60fed800800035fed301b6fe2a00e1fe00;
mem[17] = 144'h00ceff46ffe5fdf4ff5500c2007bffc4fe97;
mem[18] = 144'hfff4fe00fe3500060178fdea00c3febe00b7;
mem[19] = 144'h00b90006ff7aff14ff55007afff2ffed0015;
mem[20] = 144'h012d015cfe69fdc7016e01ebff540188012f;
mem[21] = 144'h00d9ff370088004400bbfe61fed5ff070104;
mem[22] = 144'h011cfe7bfe2600eb0051ff9bff53fdf9ff13;
mem[23] = 144'hfe5f006bfefffefeffb5ff7601af008b0006;
mem[24] = 144'hfe4200c10168fdfafe03ff760192fdfcfdc7;
mem[25] = 144'hffb9ffa6fee5017600d401a901340227ff63;
mem[26] = 144'hfe0aff510148ff80fff3fe2dffbbffd20062;
mem[27] = 144'h0145feb0fef80115004ffe9c00a4feb40152;
mem[28] = 144'hfebf006b00fbff8e0172fe98012e0169fed7;
mem[29] = 144'hfe950022ff02ff60fe85017100b8ff70fe8e;
mem[30] = 144'hfe3e00430131016f01ab0042ffddffa0ff78;
mem[31] = 144'hff8ffdfdff07ffc0fef500bfffdb0144fe2b;
mem[32] = 144'hff8f016ffea9017600810026005600c3fe6f;
mem[33] = 144'hfff7003efe920166ffbb0123fe6f0154012f;
mem[34] = 144'hfe76ff26fe68ffb1ff7b0191ff1500c90115;
mem[35] = 144'h00e9011eff97ffd2ffe0fe770174feb00012;
mem[36] = 144'h0022ffdcff0c008e0105010a009100e7fff8;
mem[37] = 144'hff7aff0a0154ff7dfe79004b006d01cbfee9;
mem[38] = 144'hff5cfe07006cff38ff98fe3801cbfeaa00f0;
mem[39] = 144'h00c8012a00f7007501ddfeee002dff4afe7f;
mem[40] = 144'h003bfeb00101feed01c601bcff1affb4fef5;
mem[41] = 144'hff95ff74fedcfe9e00d5fe6300da0004ff10;
mem[42] = 144'hfe34feda00a4fe94feeeff0fff1301de0042;
mem[43] = 144'hff6c0119013300500177016b0024ffbdff1c;
mem[44] = 144'h0100011f00e4ff6101580055ff93000aff67;
mem[45] = 144'hfe8701c1001eff36fe35fe53004c0169ff78;
mem[46] = 144'h0080ff8e01d2ff7a00f6017f007b013601ca;
mem[47] = 144'hffd8ff21fece00cbfe4601a3fe16009dfe3d;
mem[48] = 144'hfe1600ac000eff500011fe20fde00009fef9;
mem[49] = 144'hfe090079fe86ff9c002401030000ff32fd5a;
mem[50] = 144'hffc5fecdfde6ffb4fe65ff95ffb000ed00b2;
mem[51] = 144'hfe4900b9fe2c00ceff500104006afff7ffa0;
mem[52] = 144'hfe620024fd570000ffbdfdf7feffffd1fd5d;
mem[53] = 144'hfe47ff86ff9d01a001cffe5a006a007b00a9;
mem[54] = 144'hff34008aff1c0045fe94ff45fd5fff06febe;
mem[55] = 144'h00f9fe50fe58fe89fe7dff01fe5d0068fda7;
mem[56] = 144'hfda8fe88ffbe001afe32fd6e0007fd7cfd88;
mem[57] = 144'hfe41ff01003dfe84ffaafe3dfe16000e0049;
mem[58] = 144'h00dbfe52ffdb0067fef50099ff8800f0fffd;
mem[59] = 144'hfe89fe53ff9900effd89ffdafebaff4f0004;
mem[60] = 144'hfe2dff16004bfe9a0073ffc6ff04fd85ff98;
mem[61] = 144'hfedbfe7aff78fe24ffd3fdb8005efd60fe76;
mem[62] = 144'hfed0ffc7fe550064ff63ff23009aff0efdb7;
mem[63] = 144'h004fff29fe2efed1fe8f00c8ffd3fddcfe5b;
mem[64] = 144'hfbfefd53fbcffe38fccefe2cfc08feeffff7;
mem[65] = 144'hffe2fe8902fd02a201cc020b012c02c202de;
mem[66] = 144'h010402c1041304ae045f020eff0a0303fd34;
mem[67] = 144'hfc70ff23fc56fe4ffc3e019afde0ffd00010;
mem[68] = 144'hff9eff16feb800f4fc54fe53fc14ff1900ef;
mem[69] = 144'hfe8101ff0014ff7afffcfefbff83ffde0111;
mem[70] = 144'hfcb3febd00a3fe2101f40408fc03000d0204;
mem[71] = 144'hfe55fddcfd33fe96fd6f001efe8efd23026c;
mem[72] = 144'hfea4fff0ffdd030902de0341fee800c9ff8a;
mem[73] = 144'hfd81fec4007b025701250176ff4aff7f02fb;
mem[74] = 144'hff1900e1fbd8fd0c01ebfe3bff4500500410;
mem[75] = 144'h0174fe4efce9fb78ffabfdad00e6fe6b038c;
mem[76] = 144'hffddfe13fe5d002b01520020ffb500f80289;
mem[77] = 144'h01aeffb2f96df792f1aefa5dfb61f5a1fbba;
mem[78] = 144'hfe27ff84fe6bff47021403b1fff3ff460184;
mem[79] = 144'hfdf2fcf0ff8afea6ff5f002efdd101150185;
mem[80] = 144'h017cfe29fdfe01400037fe7500d2013b0020;
mem[81] = 144'hff92fefbffcb00300044fefafed8013afe92;
mem[82] = 144'hff9b012ffe01010300dc01fdfe3e00340017;
mem[83] = 144'hfefffe1a013bfe6301aafe3600bffde5fe84;
mem[84] = 144'h0068fe76ff270064fddbfdfbfe21ff950113;
mem[85] = 144'h008d005800ad01cd002b00660157007500a7;
mem[86] = 144'hff71003bfe100145005800a6ffa7ffd101f0;
mem[87] = 144'hff8b0000fe2eff5c01c100350072007801c0;
mem[88] = 144'h0005fe43fecb00ba00fe00000097ff39fead;
mem[89] = 144'hff520050ffbe00fc00d80180fe1bff3e011b;
mem[90] = 144'h00e3fe9a0016004dfdfaff930132ffbc00f1;
mem[91] = 144'h000b001ffe7eff62fe74fe3101a6006d0041;
mem[92] = 144'hff38ffd60088007bff07009bfdbdfea7fef3;
mem[93] = 144'h003cff0cfe52fe8a014900d40234fe7c0099;
mem[94] = 144'hfeab01a7fee8007e0073fff1ff28ff1bfe20;
mem[95] = 144'hfec50163011400d400410092ff61fe94fe62;
mem[96] = 144'hfc9b02d102570212030e0287fb2b0172ff1d;
mem[97] = 144'hff3501a3004300d30170033d006d01a1002f;
mem[98] = 144'hfed0ff98ff86fd49ff02038d01c3fda00081;
mem[99] = 144'h00e80173041c032701ac01a4fe2002f20011;
mem[100] = 144'hfda3001501cb03ad028a019bfc8600b3fec1;
mem[101] = 144'h02b3019200c2009fff860158008b00ff011e;
mem[102] = 144'hfcf7000b031a036e008c019afe440120004c;
mem[103] = 144'hffb8fe2f023c015b01740191fbf5ffe90210;
mem[104] = 144'hfe0bffc400c50075008c058300baff66ffb0;
mem[105] = 144'hfd9a013d019f0258031201f9fefa0193fed6;
mem[106] = 144'hff42fea5fe28fd09fe24011f03ec078b0bca;
mem[107] = 144'h021100ce02680052045c0043000104f40387;
mem[108] = 144'hff8e00bb02e9001c0006fdf0031800e60188;
mem[109] = 144'h0219fef8fa13029306b0fed9fbeef970fd37;
mem[110] = 144'hfec4013c00f402c800f103ddff3901f10259;
mem[111] = 144'hfc6aff37024b02af01740280ffcb01b30078;
mem[112] = 144'h0132012dff4f0110ff73ff68ff92ff3c0038;
mem[113] = 144'h00a9ff76fe55ff63ffecff92fea3fff70020;
mem[114] = 144'hfea9ff2afe0dfeb4fe9fff81012b007300fa;
mem[115] = 144'h0166ff8dfe77008afea00167fe3fff900144;
mem[116] = 144'hfde8010400370113ffdc00800064fef500c1;
mem[117] = 144'hff60ffd3fe4500cdffb0fed8ff410135015c;
mem[118] = 144'h01cffff900a9fee5ff35fdf900a9fed1000b;
mem[119] = 144'hff9aff9c0104feb9ff1bfed1fe32fe8effaf;
mem[120] = 144'hfe9cffe8ff79ffabff74012f0024ff3cfe78;
mem[121] = 144'hfeb3004b000afe9201720066ff590096ffc9;
mem[122] = 144'hfec0013cff0300080065fe3f008400f800b2;
mem[123] = 144'hff370061017efe4bff0000eaff69ff1afe85;
mem[124] = 144'h002a003cfe28016b00a00076fe25ff0fff4e;
mem[125] = 144'hfff0ff8cfe38013d00be01340108febfff31;
mem[126] = 144'h008cfe250094ff27ffb4fef2fe5c00c7009f;
mem[127] = 144'hfe85fdfe009000a8ff140129ff8400dd008c;
mem[128] = 144'h019d00f3fd10ffc0ff6602ed0245019afe74;
mem[129] = 144'h034d02e0fe85ff92020802ca02e10161fff9;
mem[130] = 144'h022c013300810174ffcb042ffdacfd8b01e4;
mem[131] = 144'h0017fe43ff24fe56022c014c02d0ff73fe96;
mem[132] = 144'h032e016c00a4ff3a012e00a402c2026a0028;
mem[133] = 144'h00db010cffdf01f0ffa0fe0f0072ffa700a8;
mem[134] = 144'h01bb00e3fe88ff1f009804b103eb003afe1e;
mem[135] = 144'h0199000b007bff6afe5f02190165fea3006e;
mem[136] = 144'h05cb0473ff5bfd630164049a027600530309;
mem[137] = 144'h03ad01ecfe6ffdf2ff200186027201f20126;
mem[138] = 144'hfe1402a00140fe24027a00ebffa400a305a6;
mem[139] = 144'hfe93ff9f009d00f30056fe8fffba008003fb;
mem[140] = 144'h010d007dfeb5017005ac0257000d0005022b;
mem[141] = 144'hff51fdaefb6e0188ffa8fff1010cff80fb7e;
mem[142] = 144'h017d0070fffbff4e0083032a0193ff0fff4d;
mem[143] = 144'h031c007001600067feff047002b60203003d;
mem[144] = 144'h026c00bb03b2fffffdaafbe3040401de01ff;
mem[145] = 144'h02ce0378027600820140fd6f0038009eff9e;
mem[146] = 144'h015001d70397008101b60142ffaf00b60097;
mem[147] = 144'hffeafff8fff5fdc4faebfede02ec02bc005f;
mem[148] = 144'hffd8012001c9021b0069fae1056001cd035b;
mem[149] = 144'h00710257ffde00d200bb02bd01d8026e011f;
mem[150] = 144'h03ce0239028902860150008d0322ff9201d5;
mem[151] = 144'hfec6ff18fd5f00bffe03ff57042701310128;
mem[152] = 144'h03920585047f02c90123fe980143009702a7;
mem[153] = 144'h01d8026702ab0288019ffdf403fb02780148;
mem[154] = 144'h00d4fc6bfee204ef02d2000afec0f961f0a2;
mem[155] = 144'hfd89fbc1fa9efee1fc25fdba00d7f977f7ea;
mem[156] = 144'h023301dbfe3ff990fbfa00a90047fac6fad4;
mem[157] = 144'h00db016b053e0013f907fda905170fe80ab6;
mem[158] = 144'h020e0370039901c30058fd570132fe7efe9d;
mem[159] = 144'h00ab046b01d8020501cdff4203e5027d0335;
mem[160] = 144'hfec1fe2efdc6fce80078fed8fb4b00a9003e;
mem[161] = 144'hfd1effee00c000c40026ff59fc8e01ff02b4;
mem[162] = 144'h016702dc01bc01b30157ffbbfe02004d0187;
mem[163] = 144'hff060013fd6d003bfdc600ccfe10031f0125;
mem[164] = 144'h0012ff97fe0dff4b0032fdb2fe42fefa03a3;
mem[165] = 144'h003afe7d00c4025c008c0116ffbbfe7effb1;
mem[166] = 144'hfcbffddd00a7000cfeda0213fcc600f10221;
mem[167] = 144'h019dfcbffe01fdfd0034ff63ff0800940376;
mem[168] = 144'hfce9019cff4d013bff5bffd3fd9e034d01ba;
mem[169] = 144'hfd80fefe0078fdf0fff9003ffb66003c0345;
mem[170] = 144'h0386016401f6007203e3ffef029703630445;
mem[171] = 144'h02540039fd50fbe70053fe7d0311017c0684;
mem[172] = 144'h01dcfff3ff1c0258008b028301d605480265;
mem[173] = 144'h01d4013efdd3044402ef00d2fe05f9f402eb;
mem[174] = 144'hfd7e0104fce300cf0014013efbfd0332010a;
mem[175] = 144'hff30ff1d005200e6ff31010ffe6a0333017f;
mem[176] = 144'hff44ff58fe02ff45000b00eb01aa004500d5;
mem[177] = 144'hff6cfe41ffc8001d00fefe2b0160012aff5c;
mem[178] = 144'hfe1800fbffbdff18ff3fffc9fea100e600e4;
mem[179] = 144'h00cbfde50073ff8e00f5ffb8fefdffadff98;
mem[180] = 144'h016b017afec3fddfffc700b701b500d8ff8a;
mem[181] = 144'h0069fe4300210073ff8b016f006afe9700d9;
mem[182] = 144'hfe2bffe8ff1f0017fedafebd00afff65007b;
mem[183] = 144'hfeb3014f01d5feb60034fe5b0091008001dd;
mem[184] = 144'hffdbff0400deff960134ff9400b5ff8fff92;
mem[185] = 144'h01d2ff89fed0003cfe08009600f8011a0216;
mem[186] = 144'hff78fe41008f003dfe8e00cbff460090ff54;
mem[187] = 144'hfe0200bfffd6ff89ff82fe48fe29feb6fe43;
mem[188] = 144'h014cffc1013d000fffacfeffff67004f00f4;
mem[189] = 144'hffc9002c006aff93003eff9cffff003afea5;
mem[190] = 144'hff14fe4f011aff98ffadfff3ff0d01bafee6;
mem[191] = 144'hffef00fc0049fe33ff7b01010063001900d9;
mem[192] = 144'h019602dffff7ffd90169028f0234005d00af;
mem[193] = 144'h012cffc8ff3dfdd3007c0299ffef02ca00c0;
mem[194] = 144'hffe5ffd3fec9fc8ffff200abff17ffa4fd93;
mem[195] = 144'h02590027fe5a030d02d303ee026e0017fdc2;
mem[196] = 144'hff08013efe22feb00168041100df01aaff25;
mem[197] = 144'h01530090018400eafdd200d5013dfe2cff72;
mem[198] = 144'h00c7007ffebdfedb0055029c025500000058;
mem[199] = 144'hfdc6028e0202ffec02880227011dff0aff85;
mem[200] = 144'h0277001dfe72fded03160557fff20293ff43;
mem[201] = 144'h02cf00b8ffe0ff35006e02f701430197fe92;
mem[202] = 144'hfe7bfd49ff2ffbb1ff79010efdd6fd31069c;
mem[203] = 144'hfff2ff3002ad026b007e0076fe85034803f1;
mem[204] = 144'h02d8ffcb007d03910421ffd6fed50192001b;
mem[205] = 144'hfe27fc04fba4fbc0fc05fcad01ce00a8fa6a;
mem[206] = 144'h011d030dfdcf00b8008201a6036902a200b3;
mem[207] = 144'h017e004600c9ffd5020c035003740080ff93;
mem[208] = 144'h00b1fa92fd79fa8afd0f0086029f010b00c6;
mem[209] = 144'h008a0042ff6bfeb700f102d1002eff47032a;
mem[210] = 144'h01a901340573013a02a502bf004b01fefd13;
mem[211] = 144'hfe64fb3cfc42fd70032104f400d2ffaf0312;
mem[212] = 144'h040bffe7ff75fd56fe2aff25020c00bd0122;
mem[213] = 144'h00cafe5801bdff02fdbbfdc100a7fe3d0110;
mem[214] = 144'h0035fc96ff90fdc70068015c0295fe8f018a;
mem[215] = 144'h00e90039fde3ff8efd51ff5101f600080342;
mem[216] = 144'h02ff017301b7004e00de0185ff22001f0057;
mem[217] = 144'h0302004c00e1fcb8fe9bffe5012701d002ce;
mem[218] = 144'hff8b00cf01df040fff1c027c021affc80135;
mem[219] = 144'h000200000193ff80ff65006f017d01cd0252;
mem[220] = 144'h00b0010600bc011e051103e8ff6701ef0071;
mem[221] = 144'h01f1ff76fb93f90cfb23000704e103450064;
mem[222] = 144'h010eff3e0165ffd8ff20028b0122ff6aff2a;
mem[223] = 144'h0182fe3d00d0fcb5ff38031f00fc007201ec;
mem[224] = 144'hfe7801c4023e00d4fc62f9ba00fa044e05cd;
mem[225] = 144'hff2c039a0452049bfefafc8b02bc0253007e;
mem[226] = 144'h004000e003ce0383041d007701f5fde2ffdb;
mem[227] = 144'hfd860260003ffdc4fac1fdc001180476ffd5;
mem[228] = 144'hfe69fe6503040326ff68fe2300b7018a00ec;
mem[229] = 144'h0155000bfdf8ffb4ffd502d1fffb024dff18;
mem[230] = 144'hfd0903020560029a0320fd12ff7d04b90362;
mem[231] = 144'h004efd6afc4bfd82fd75fc59fd47025000ac;
mem[232] = 144'hff93036106c6042801f0fc3b02c703c9006a;
mem[233] = 144'hfcf603e2038d046902ca00000048030902ce;
mem[234] = 144'h00a0fd50fc2bfe41000f00e1002dfb4cf221;
mem[235] = 144'hfecdfcf9f5f2fa0efd3afc95fd92f97cfa7a;
mem[236] = 144'hff49033afe90fc9bf4c000050338fed7fb49;
mem[237] = 144'hffa901a902d7010bfaa9fe2e00450bcf0fdc;
mem[238] = 144'hfd66007902ef050c02a3fe43fe790260013b;
mem[239] = 144'hfd3801a901ef04980010fee6fe4802bb01ac;
mem[240] = 144'hfc24fd5bfdafffd3006f0230fb4a001b0093;
mem[241] = 144'hfd62fd280007006f032dfffffdc601a10117;
mem[242] = 144'h011bffefffe401c0002a00f7ffc1fed503ee;
mem[243] = 144'h017300b0018801ad04e8034cff1e022f056f;
mem[244] = 144'h00a3fecffc27001f023402e8fce6fd21ff7c;
mem[245] = 144'hff79ff61016400d00214ff6b00ca01af0164;
mem[246] = 144'hfe1efde3fde10127014100c9fe0afff8006b;
mem[247] = 144'h026e00b0ffc4024d01590362fbb0fc8701b2;
mem[248] = 144'hfc17fd4701ad0375003200ce006301a30068;
mem[249] = 144'hfc78fb4cfea8030a00be03e8fcdb0063ff28;
mem[250] = 144'h03ab0509067dfda8026cff9b067c09020ce4;
mem[251] = 144'h03a004a4042402600361022803ad038504d0;
mem[252] = 144'h0128014305e8061703ecfefb02b304580982;
mem[253] = 144'h030700d4f8b100b005a305e6f9feeedef604;
mem[254] = 144'hfd34fe00ffb60178047d0258fee1fe490182;
mem[255] = 144'h0125fc90ff6500a8020703dbfe0cffc701a5;
mem[256] = 144'h03cc0239024c04ed024802350215011b00dc;
mem[257] = 144'h018001df0121016bfebcfff601abfdbf00a6;
mem[258] = 144'h0009ff2ffee5fd11ff750098020cfd7b02ee;
mem[259] = 144'h012e036904b80207025cfe8a003a01a100ea;
mem[260] = 144'h00bb00cd01230294030d01dbffe70008005b;
mem[261] = 144'h002100640130ffcb015bff4001d4ffe20263;
mem[262] = 144'h002c027c0189030efefeff1400d401d10068;
mem[263] = 144'h00b2025700c403110379ff76022bff02ff90;
mem[264] = 144'h029201f1fe76ff7d010d0347025b00a50191;
mem[265] = 144'h01b3ffc2011800c0001e01610145ffc50009;
mem[266] = 144'h01a900f00367fe92008f016f0176021efeb3;
mem[267] = 144'h024a0222019800e6026101deff930297009e;
mem[268] = 144'h00360172034402a6ff6400c001bbfff70286;
mem[269] = 144'h0105febcff2b05c70a320656fdabfc62fc28;
mem[270] = 144'h02d7016b01a20217007201f802670208fec8;
mem[271] = 144'h003cffe2ff320189031c01a401abffb100b0;
mem[272] = 144'hfd8901b502f203900249ff32fdb000760146;
mem[273] = 144'hfec9fe1001140135fd9bfd13002c02ea016f;
mem[274] = 144'hfe5fffa5fde4ff0cfdaf001702e0ff140317;
mem[275] = 144'hfdaa01f8032003c0003cfee3fe3602fc0117;
mem[276] = 144'hfdda0030004d02c1038002c5fb8a00a4fefe;
mem[277] = 144'h01c501cdffc50097030c0073005202c10220;
mem[278] = 144'hfdfb0083ff00022f0143fd7cfe8e018402d6;
mem[279] = 144'h0008ffe7fe0602e901e30198fcbafe3f0036;
mem[280] = 144'hfc720013fec201a4ff6ffe61001e03fdfe1d;
mem[281] = 144'hfa8f0038008d020f00e9fe57fd7d0035fec9;
mem[282] = 144'h002100b302e9fd7ffecd0036027205e70631;
mem[283] = 144'h008e030cffb00076052a01390194029803e4;
mem[284] = 144'h0104036e02d900ebfdbdfd5001e902a000fb;
mem[285] = 144'hff71fd78fe4f05f90b6a05a1fb90f85402b8;
mem[286] = 144'hfdcf00f601b80344ff5afe8d00050378020a;
mem[287] = 144'hfe1a007c01b701a1013cff7efbc8ff25ff5c;
mem[288] = 144'hfea0fde1ff9a00a201ad02b0ff9e00900111;
mem[289] = 144'hff790002012b0294027b0369fdec0259fd7e;
mem[290] = 144'hfffc00210165049b0108050700b000c7fb6e;
mem[291] = 144'h000dfd5f021c003800fc0257fe2effa7021d;
mem[292] = 144'hff7eff0e00a301d7000efe9effbafded016f;
mem[293] = 144'hfe74ff00ff34ff3e0103fe3d006d01e100cd;
mem[294] = 144'hff80fd47008c007c011f0285ffbcfffc02fb;
mem[295] = 144'h0163ff5a018b010c008101d9006300c00298;
mem[296] = 144'h0076ff62019a045602a306020059002cff6e;
mem[297] = 144'hff6d003201ef01cd008c021affd6ff9f0083;
mem[298] = 144'hffbb000dfb25fadc02550155018d012a056a;
mem[299] = 144'h0131fee5ff90feb70272fffb02bf01790483;
mem[300] = 144'h004f01d10159fe940154007dfeea022b01e4;
mem[301] = 144'h00cdfdd6fb660046fae9fca7fde6f94afdf0;
mem[302] = 144'h019dffd60408025701150273ff7cffaa0137;
mem[303] = 144'hfecbfe1701ce034800640138fdb1ff71021d;
mem[304] = 144'hffaa000d0045fe8e00870078fffd007d007b;
mem[305] = 144'hfe15ff81fdd8fe1500940012ffc500a30059;
mem[306] = 144'hfe4a0111ff09ff35010d0024fe2900290104;
mem[307] = 144'hfdcd002aff4700a2ff2d0072ffc3ff5afed4;
mem[308] = 144'hffe0fe9dffc7ff46ff4ffe69003fff700018;
mem[309] = 144'h011a01770148004b00eb00e10153fe93ff68;
mem[310] = 144'hff49fedffea8fdb1006200d300a5fe690134;
mem[311] = 144'hfea9ff65ff37006000a6fe4100fc0034001b;
mem[312] = 144'h0119ff6b0032ff23ff21ff0a002900f10160;
mem[313] = 144'h0020fde9feee00ed014b00d300f80097fe92;
mem[314] = 144'hfe36fe2afea60097ffaafe1effbdfef800be;
mem[315] = 144'h0023005cffb8febeff2100130140007dfdd2;
mem[316] = 144'h0087fe49ff5e00200110fe140059fe3b00ad;
mem[317] = 144'hfe3b001a009eff83ffa70140ff5bff63fef6;
mem[318] = 144'h00f5014e010b005d00f3fdfcfec100a7fed8;
mem[319] = 144'hfecfff62feb0ffbdfe9100bf014ffec6ff4c;
mem[320] = 144'h03d7fd0afebffe8a002f01fa00effbf9fcc4;
mem[321] = 144'h0380fd84fdcffeb5001bfe9bfd0cfec001be;
mem[322] = 144'h019800f002bbff9a0154fef501200149fecc;
mem[323] = 144'h01f3fc4400ba0236045103dffddbfd7003a1;
mem[324] = 144'h03de0055fcecfec0fe05fea801d9feb8feb6;
mem[325] = 144'hfeb4ff00fde0ff22ffc5ff84ff38fdbeffae;
mem[326] = 144'h0326fdffff6e00160110fdd9fee4fb72fdb5;
mem[327] = 144'h030000b8008a00bffec9ffed031100a0fe97;
mem[328] = 144'h005bfd75fe16004a0002fda6fd28fd0b007c;
mem[329] = 144'h01adfd13fd91ff00005700a1ffccfb85ffa9;
mem[330] = 144'h028700830551079300e9018000cf02ed0190;
mem[331] = 144'h00bf0307037a03b0015e023600ef0344ffdf;
mem[332] = 144'h010effc503df05fc05d2027bfd9d00ed0461;
mem[333] = 144'h02b303d7fdf8f9f1fdc6023f024d0189fbc4;
mem[334] = 144'h047afd93fe42018fff37fe6400b2fe29fdf6;
mem[335] = 144'h0449febdfc4e0043010c0022ff39fdf9fdbc;
mem[336] = 144'h01d100bafea3fdcf047e06f001f4015afe13;
mem[337] = 144'h0236017cff3ffef800f7049f00e8008d0026;
mem[338] = 144'h017d03d9ff1bff4dfe3f0209013ffd5803aa;
mem[339] = 144'h01a0fdbd011a03b704930504016901520023;
mem[340] = 144'h00fe00abff2dff42024402c30177025201af;
mem[341] = 144'h007100c1014bfdf1005afdb40148fe050040;
mem[342] = 144'hfff5013afdfeff5200f80382021301c9ffea;
mem[343] = 144'h0068003f0134001101b502f1fdc3fe7f007d;
mem[344] = 144'h020e02eaff4cfe7700be0695ffad00ef01c9;
mem[345] = 144'h03850285ff7cfcb6ff8905e4ff7402eb00f5;
mem[346] = 144'hffef02950537fcfdfe31ff88ff2e01ad0c8e;
mem[347] = 144'hfee100a8062f026900ea02190253038d09f8;
mem[348] = 144'h0117ffbbffcd02b0072b017a007e0345034c;
mem[349] = 144'hfe24f978f87effbd062e01a60011f7c8f917;
mem[350] = 144'h0267023ffe77fd98024b05b702a9022a0048;
mem[351] = 144'hfff600e0001cff88ff3f02c000a401a00024;
mem[352] = 144'hff42006afe18001cfef60087fe1bfe95fde7;
mem[353] = 144'h016c01bdfd26fef4ff38ffadfaf4fcdcff45;
mem[354] = 144'hff3000870009ffba01880217fd1f01fb0362;
mem[355] = 144'h012d00dbff0ffde4fd9b0004fd6ffdf4fe9e;
mem[356] = 144'hff2700a8008cff4d000400460104fd69ff84;
mem[357] = 144'h0052fff101860232017ffff10060ff2b017a;
mem[358] = 144'h01b80112ffaefe4300930156febffb7afce4;
mem[359] = 144'hffe9fff10289fd28ff87ffd401e90021ff92;
mem[360] = 144'hff21fdecfd58fea6015c0052fc80fcb1ff86;
mem[361] = 144'h018401d9fcf9fe62ff9a02b7fb75fda2ffd3;
mem[362] = 144'hffe101af03ef003a00bd01fe02e605b70406;
mem[363] = 144'h00d301df01f80047001a01740382004f022a;
mem[364] = 144'h012a00e1fef502ab06910134fdbd0162ff05;
mem[365] = 144'h009f033d0637ffe6f8d0fe7c01fc039b017b;
mem[366] = 144'h01000148fe66fe22fe6a00cbfd44fd96fd0e;
mem[367] = 144'hfea200350021ff02fe8cff6efcc6ff26ff1a;
mem[368] = 144'hfebd0006fe86ff020166014d01b2ffe500d5;
mem[369] = 144'hfe5cff83feda0057ff03fe31ff6f01980089;
mem[370] = 144'hff72ffca0187ff730075002d01bf003afe6c;
mem[371] = 144'hff2bff4d0095ffdb009afedc0187ff1cff31;
mem[372] = 144'h0174fe8f010ffe11fed7fe2c01dd006e005a;
mem[373] = 144'hfe33fff80006ffcd00e7ffdb0176005dfef9;
mem[374] = 144'hffe10142fe22013aff8100cf004200d2ff6f;
mem[375] = 144'h010bffd70101ffef0059006001140172ffc2;
mem[376] = 144'h005a0042ff7b0095ff93008aff7fffd2ff2d;
mem[377] = 144'hfe80008400adfe25ff4cfe990139fe1f00fe;
mem[378] = 144'h00a9018dfe65ffb0011e00bafe69009bfee0;
mem[379] = 144'hff7800cefe5afe0cfe13fef4ff4dff71ff29;
mem[380] = 144'h0131ffaafdcc0061001f0052ff4bff0dff19;
mem[381] = 144'hff88fe8f006a0110ffa2ffee005a010bffbc;
mem[382] = 144'hff61ff8b000a00fa000b019cff2601b7018a;
mem[383] = 144'hfeb4ffedffcb008600a2fdf7fdf80171fe33;
mem[384] = 144'h0062fedcffb8fdeb00800073fefeff30fd6b;
mem[385] = 144'hffd4fe81ff4cfe490015ffea005900c6fe6e;
mem[386] = 144'h0067fff4ff21ffbd0036ffee007700f2ffc8;
mem[387] = 144'hfc8ffd4bfd47fdaf0108fe300040ff94ff02;
mem[388] = 144'h0051fe0cfe14fe3bff37001afef10074fe11;
mem[389] = 144'h00350132ff7eff0401610092ff9501a10118;
mem[390] = 144'hfd19fe62fd4dfcf7fe9000d3ff1eff280120;
mem[391] = 144'h0018fca7fd1b0044fe8cfe42fe76ffaa0046;
mem[392] = 144'hfea6ffd9fddcfe8c007cfe9e00af0049ffdb;
mem[393] = 144'hfd17fccffe6500170010ff68fe3cfebdfd99;
mem[394] = 144'hff9001480113fef5fd5600f5fdfd004300aa;
mem[395] = 144'h000cff70ffb8ff79fea5fdbffe45fdddfef6;
mem[396] = 144'h00dcfee7fe1afe94013b009cfe7cfef7fea0;
mem[397] = 144'hfe5dfe680041005f0108fdf9ff10fdaf001c;
mem[398] = 144'hff12fef3fe7cffbf0018fe67fff1fe13fe4d;
mem[399] = 144'h0062fe74fd47fd26fe15fdfb0030fecafecb;
mem[400] = 144'hfe55fd89faf7fe1ffd7efd5afe0cfceffd8e;
mem[401] = 144'hffb4017cfddbfd3fffe7fe1bfde4fd190140;
mem[402] = 144'h0084031a02350163ff96fee1fde00255013c;
mem[403] = 144'hff29fd63fa7afac3fcd900c5fd890011ff89;
mem[404] = 144'h0057ff430137fdeffc5ffc6501c4fd600342;
mem[405] = 144'h002ffd9b005afdfafd14fd60fd59fd470068;
mem[406] = 144'hfe6a000cfda3fdb7fcadfdc0fef5fe80fcd5;
mem[407] = 144'h00f300f6fe3ffd43fcfcfc260021fd9d01b3;
mem[408] = 144'h00a0ff90ff58ff9efc02fd0efce7ff0affd2;
mem[409] = 144'hff5400aeffa0fe75fd6dfc87fdf6fee2ff1c;
mem[410] = 144'h0154017400ae046b02faff0d004f02aefe7d;
mem[411] = 144'hffc2ff0b00eeff8b0072fce80135ffd0008d;
mem[412] = 144'hff75ff56fea6fe8902f50339fdaa01deff4a;
mem[413] = 144'h014b0183019ffbf9fbe8feb4040904ed024e;
mem[414] = 144'h0064fd920036fd73fd1dffe3fda3fd16ffe1;
mem[415] = 144'hff13fff4fd98fe66ff17ff2dfe9cfdb40154;
mem[416] = 144'hfde4ff10fdb400a3ff39ff87fb88fe12fe36;
mem[417] = 144'hfcdcfe6dfdf9fe00007eff25009aff75ff35;
mem[418] = 144'hfe56ff8bfd6dff0dfd57fdfbfe90fe4cfdc6;
mem[419] = 144'hfef7ff22fea3fd97ff2dfdbafc540189fedf;
mem[420] = 144'hff41fbaffebc020401a5ff0cfc9affa900ab;
mem[421] = 144'h0052ff7d00f2009a017201c100eaffedff15;
mem[422] = 144'hfba3ff37feb3fe5dfec2ffbafe3cff71fef8;
mem[423] = 144'hfe7cfcc0ffc20162ff23fed1ff46fe4fffb1;
mem[424] = 144'hfd0bffceffc8fe96fded0056fe3d0026fbf0;
mem[425] = 144'hfd1efc9c0051ffd80041fe58fffbfec3fef2;
mem[426] = 144'hfc2cff77fd2afc79fdf6fd26ff12ff3efec9;
mem[427] = 144'hfcfefd05fb71fbad00c2fd62ff10fd6ffed0;
mem[428] = 144'hfc65fedafd85ff0ffd35fd67007dff90fbfe;
mem[429] = 144'hff90fe4400900014ffa6fec1fe29febeff3f;
mem[430] = 144'hfe20fe80ff16007d0057fe00ff11ff2cfe44;
mem[431] = 144'hfe0afd62feb8ffff00a3fd16fcc2fe5ffea9;
mem[432] = 144'hfec0fee3fefb0174002cfde7fe1cfdfe0155;
mem[433] = 144'hfe6effe801280160fe85010c01ce00f300cc;
mem[434] = 144'h00310058fe22000cfe9900eafe30ffb8ffd9;
mem[435] = 144'h004cff38020d002800790074fdad013bff24;
mem[436] = 144'h00a001380089fde5ff4dfe59fffcffd900ce;
mem[437] = 144'hff87001701b800f30008000e010f014001b0;
mem[438] = 144'hff46fe8e006a011aff71ff33fe08fdb7ff52;
mem[439] = 144'h00d901dd013e00f7ffdc0143003d0029ffbb;
mem[440] = 144'hff6e00e9fe41ff51fe6500e3ff7a00fafdb8;
mem[441] = 144'hfdf6ffb8fe10ff3efe55010cfddf00060144;
mem[442] = 144'hffd9006f0045ff2aff70011e00e60233ff89;
mem[443] = 144'hff88fecbfe810223fef90007fefb01040217;
mem[444] = 144'hfded002f00eaffe1ff42fe28fe52fe5aff3c;
mem[445] = 144'hfeb4fdbf01380102fe050176fe9afdafffea;
mem[446] = 144'h019400affec10181010cfe4800f80021feb3;
mem[447] = 144'h007efe2efe22fe6cffd1fec10064006c00af;
mem[448] = 144'h01b000fe0179ff7600acfefdfefdff350077;
mem[449] = 144'hffdf01a000f500420072fe8900c701abff9a;
mem[450] = 144'h00a5ffaf006efdc9ff4a00780123004cff4e;
mem[451] = 144'hfea9ff84009cfea2ffbb002600fb0031fe44;
mem[452] = 144'h00eafe510148fefb006aff2effdc0066ff9c;
mem[453] = 144'h0077ffe2001efff40116ffec00d0015300b1;
mem[454] = 144'hff5effa4010dffa800af0094fe96ffd1ff0e;
mem[455] = 144'hfeff01ab014bff57018700fffe6500c6fef8;
mem[456] = 144'h003c00e2fe6801400095fdc8fe4a0108fe3c;
mem[457] = 144'h014dffeefdeafe71fe8f00c9feb8009bffe3;
mem[458] = 144'hfe6affae0154fde3015fffd7014c022cfec6;
mem[459] = 144'hffecfe29001dfdffff5b000bff40009b0150;
mem[460] = 144'hff4cfeeeff8efdc4fe22fe4dffff0068fe00;
mem[461] = 144'h00fafefffe5cffe100f7febb003f022fff68;
mem[462] = 144'hffdcffc60187002cff4800140094feb801cf;
mem[463] = 144'hfecfff19010400220124ff32ffa5ff32fe5c;
mem[464] = 144'h003904230095030bfd7eff4503fe02a202fe;
mem[465] = 144'h01a1029c01dc0017fdbefe0701fe00760187;
mem[466] = 144'hff4b002e0062ffd1ffd5fd58008fff66fffe;
mem[467] = 144'h02640286febb008ffd9afee5038c0141fe62;
mem[468] = 144'h006f0214ffb3011d000d00fe0272044e027e;
mem[469] = 144'hff160183ff2dfedcfd7001e4ff540000ff12;
mem[470] = 144'h02a2042001cd0121ff88fee5026f0204fefb;
mem[471] = 144'h007fffb1001b003cfe23ff9700de03330196;
mem[472] = 144'h039600d4026400d2fdbdfd55026601e5ff9a;
mem[473] = 144'h01dd046602cf0021fe73ff9100d102cf0344;
mem[474] = 144'hfd2afd8eff0dfd6b0106fe75fd97fba9fb42;
mem[475] = 144'hfef4fc4aff34013b0113002fff37005bff9c;
mem[476] = 144'h02a9002a0023ff6cf942fda6001b0060fabb;
mem[477] = 144'h000cff5f00f4012500540262036d03f0061b;
mem[478] = 144'h0084033eff9f01a4fd49fcfbff9300c8ffe0;
mem[479] = 144'h00e603b3017b02a3fed6ffdc00720195029e;
mem[480] = 144'h000800ed02e103fcff5dff0f00c2004700df;
mem[481] = 144'hfe7c012c02870224005bfe09002202daffe9;
mem[482] = 144'hffcf01dc0101022f00e2fee2024e0367fb77;
mem[483] = 144'h000d0204043affb701fcfff302190054016e;
mem[484] = 144'h0140013f020201b801ab0058021e041a0078;
mem[485] = 144'h003a004b000ffe68ffc1fe3501c900d3005d;
mem[486] = 144'hffeb025a01fb0283ff19ffb80047fedaffe5;
mem[487] = 144'h024202c200ec029a013702d70198025afd1b;
mem[488] = 144'h01ac000b02de01030101fca201cc00ea014b;
mem[489] = 144'hfe9effb101ae008002fcff7d005201e1fee5;
mem[490] = 144'hfe83feedfb7b01c6ffe60008feadfe860394;
mem[491] = 144'h0062ffa2003a0394ff78033cfe7f024afe81;
mem[492] = 144'h002f0245025afef5023b0105ffb702b0fb95;
mem[493] = 144'h008c0048ff82fb79fa94ffbe00190487013f;
mem[494] = 144'hffc8025603740325ffebfcd7fef302550023;
mem[495] = 144'h017e007a027f02c000fb013902c30278012a;
mem[496] = 144'hffddfe15007d011ffeb0002bfe4e0048fdbe;
mem[497] = 144'h006cff97fdcf018d0077fdfb0153fe3000fa;
mem[498] = 144'h0031fff500bc015e0103fdbcfdc9ff2bffad;
mem[499] = 144'h013cfea6fdb000530011fee7fdc2fdc1fe3b;
mem[500] = 144'h0067fe890135ff3300b80186ff4bfdc2ff3d;
mem[501] = 144'h01bd0006fe6dff6a0022fefb00edff6301b9;
mem[502] = 144'hfe4600e5ffb8ffd2fdf1ff6dffbbff7c0069;
mem[503] = 144'h00bd0121fef8ff61fe09fdb3feef0190fee8;
mem[504] = 144'h0036000a010700c9fec4011100d8feb8000f;
mem[505] = 144'hffe8ffd20064fe23fe8800e4010dfd97014d;
mem[506] = 144'h005dfea6021afe43ff2400c1fe55fe49ffcf;
mem[507] = 144'h00dbfee300eaff0f003d0150fe82ffcd021d;
mem[508] = 144'h0096012c00e10086ff89ffa900dcfe4cfe18;
mem[509] = 144'h0045fef1fdd800f60003fed6fde8002b00cd;
mem[510] = 144'h00ea019b0037fe67015801c901550076fec5;
mem[511] = 144'h007affcdfde70003fecdff43fdc500ffffba;
mem[512] = 144'h0074004d00f6ff10fa4cfb9fffe7040c01c0;
mem[513] = 144'h009b0126028afe25fbbcfcd801f505cf01e9;
mem[514] = 144'hff6000630417021ffd6cfe6f03e801a30170;
mem[515] = 144'h017400790040fd8ffc9ffd6d01f8028600fb;
mem[516] = 144'hff6b02340184fe77fd75fd40010601690330;
mem[517] = 144'h018b0014fe5bff6aff1cfe4100ee0116fee5;
mem[518] = 144'hfe2b02aa0341fffdfdb3f9e4034f01950317;
mem[519] = 144'hfed8ff660131ff72fdf7fca6000e00d100bd;
mem[520] = 144'hfe7002cc02fe0086fa70f88b03f9051402fa;
mem[521] = 144'h00f9033b0357fe58fa7ffc94013902ae040a;
mem[522] = 144'hff6f0128fedb0743021a0057ff73fc9cf69f;
mem[523] = 144'hff4dff6efd5b0354fd86fcb6fdc7ff2dfee5;
mem[524] = 144'h028802c600c2fa64ffd20298016a0408fd7e;
mem[525] = 144'h023a01cb00ddfb88fcf501eb01b2017d0248;
mem[526] = 144'hfefb0227027dfdc7fb84fc0d00e504840279;
mem[527] = 144'h0055009f018fff29fe43fd74024d030102a9;
mem[528] = 144'h0072fe3aff13fecb0034ff33fca4020a03f4;
mem[529] = 144'hffbbff5a02bb01b1fff202f60137024e0158;
mem[530] = 144'h0185024201b5040d037004e300050267fc04;
mem[531] = 144'hfec200f3fe4cff5efd2500beff3905470056;
mem[532] = 144'h00f3fed001090129fe6efeccfd0502610214;
mem[533] = 144'hff0cff54febfff9d0072ff71005e003d01b6;
mem[534] = 144'hfca5ffcf034300cb02e602e0feed03570468;
mem[535] = 144'h01660020ff7eff6efe27ffaafe99ffc503b2;
mem[536] = 144'hfe3a027504a701a400ae03eb01cc02bf0217;
mem[537] = 144'hfe3e00af0223011affe300a4fdcf021f02cb;
mem[538] = 144'h01a00136ff2bfd300270ff4401b1fd890069;
mem[539] = 144'h029d026afdf5fb1d006eff3d03fbfefd0337;
mem[540] = 144'hffa0033f01c3fc490029014b039a066400c5;
mem[541] = 144'h00b70071fe5903a3ff1efd78fe7ff3f10245;
mem[542] = 144'h0064ffe6032affe401cf04a50164051e0175;
mem[543] = 144'hffa4ff760240008701e10102fee304cc03f8;
mem[544] = 144'h015a004e00fbfecefec0fe8ffe4d0085ff0c;
mem[545] = 144'hfd9ffdd7fefcff84fe56005e0123ff300084;
mem[546] = 144'hfedf0052008e0085014e00e9ff2300efffd4;
mem[547] = 144'hfe7afe69ff17fe6efed9feccffff0031ff4f;
mem[548] = 144'h002cfe9ffe66fe47fef8fdedfe70fe060063;
mem[549] = 144'hffc9ff4c01970006009300bf0170fe410128;
mem[550] = 144'h00a3fdeffdf5012fffdafdc2fe67feecff9b;
mem[551] = 144'hfee5ff5d01120087ff3dffe5ffe700c900ee;
mem[552] = 144'hfdff0128ff2b013f0042fec00076fe2d004a;
mem[553] = 144'hff6ffe9fff91fd9ffec0014c007cfe78fda1;
mem[554] = 144'hfea0ff5fff5d010afe30006400e2feba0119;
mem[555] = 144'hff4c00e4ff0f0156fef7006bfe1ffecfff0d;
mem[556] = 144'h01490062ff5dfde1fe7effa6ff8cffc5fe6a;
mem[557] = 144'hfe24ffeffdec0069fea2fdb1fe8b0150fdf4;
mem[558] = 144'hfe1800defdeb00a1fefbfe34fefafda800ae;
mem[559] = 144'h014efe43fe4f0142ff92feec00c5fef10000;
mem[560] = 144'h0400ff3e02af00e9ffdcf8a601fb034004c1;
mem[561] = 144'h029501c00331017a01b5fce002c3febbff2c;
mem[562] = 144'hffecffb803b101b702ecff8802d2fdccfc53;
mem[563] = 144'h0012ff8c0093fe17fcf5fe0d0238ff5700d8;
mem[564] = 144'h0110011202fa01e3fea6fd3103f00128ffb8;
mem[565] = 144'hff96016d002a00d702d40200006b017f01b4;
mem[566] = 144'h023901fe021903db001cfc9002f901060283;
mem[567] = 144'hfe790012fd5501590083fe3602e7017a001a;
mem[568] = 144'h0292029302710280017af95c0116ffa30246;
mem[569] = 144'h04270029020103b0016efc08022c014e011b;
mem[570] = 144'h011afedffd0202a000be0047fe48f6e9f04c;
mem[571] = 144'hff16fe8afba5fcf9fd260034003bf974f782;
mem[572] = 144'h012300a701c1fbd1f5eb00fa00f4febefdf3;
mem[573] = 144'h005c043c01edff56fb38ffd302e507c706c0;
mem[574] = 144'h037dffe700a2034401b0fc3002aa012fff82;
mem[575] = 144'h0237ffba035802b302a4fd6b013600fb0096;
mem[576] = 144'h006f02cbffdcfdf8fcb2fbdf063a04a2029d;
mem[577] = 144'h00a601c80187005601bdfe7301c10071ffac;
mem[578] = 144'h01330019034c0203035d0088021dffd1fc21;
mem[579] = 144'hfe7b01cfff4ffccffa02fe4800770262020b;
mem[580] = 144'h00d6013b00a401cc013afab70323049e034e;
mem[581] = 144'hff7dff32fec9ffbe009a00c4015e01e0ff6e;
mem[582] = 144'h02ba024104e501030235fcbe05bd01ce00d5;
mem[583] = 144'hfd55ff88fce5fdd8fef5fe2d0173031d0136;
mem[584] = 144'h033304b604860484025efd62049601720263;
mem[585] = 144'h0462041f038a030d01b9ff0d0557042c028a;
mem[586] = 144'hff4afeaefb95fe0e033bff15fad7f8baed2e;
mem[587] = 144'hff4af9a4fa4afbb0fd7cfebefc77f92ef828;
mem[588] = 144'h00c00230ffc3fe44f658000e012bfdfdf913;
mem[589] = 144'hfd00ff9c025bfa29f65afb8e016d09e006e4;
mem[590] = 144'h00f000e90321037eff7ffd1e04410014ffb1;
mem[591] = 144'h00190206049d03e00245ff18039e02440333;
mem[592] = 144'hfe95ff01006afff7ff2bff090015fe840145;
mem[593] = 144'hfeed001a0131ffe0fff101cbff72ffaeff62;
mem[594] = 144'hff66013aff69ff310062fecdfdeafed40227;
mem[595] = 144'hfecafe8afeb1009bfe070194feeffe1efecb;
mem[596] = 144'hffeffe540107ff14ff22ffb10054ffcdfdef;
mem[597] = 144'h01d3ff5a006a00b6ff2cfef5019bffe10068;
mem[598] = 144'h01280016fe36002bfe9eff750060016afe76;
mem[599] = 144'h01450068ffdb000a018500befe92ff43ffda;
mem[600] = 144'h009affa9012b00a6ffc40139007a016afe9a;
mem[601] = 144'h00a8ff5dffca012dfdbdffa1fdc9ff8ffe24;
mem[602] = 144'hff560045017700610103fe6a00770015009b;
mem[603] = 144'hff06ffd40103ffd3013801c8fe9cff6afe75;
mem[604] = 144'h00d40113ff340015fe75fdf50025008fff66;
mem[605] = 144'hfeadfdc2ff43013101fefff2ff99ff85ff0c;
mem[606] = 144'hfeb7fffa01df0129ffc1ffe1006f00d60183;
mem[607] = 144'h008f0065fe76ff52ff33ff2cfed6feffffbd;
mem[608] = 144'hfd6bfc9afebe00ef0036fbf7fee800a0fff7;
mem[609] = 144'h000501cb0167fed7ff0800b001390146ffe8;
mem[610] = 144'hfed4ffb90287fff40138024500d30042ffd2;
mem[611] = 144'hfe8dfeba00efff5ffd5bfc8700080361ff63;
mem[612] = 144'hff84ff0600a4ff0501e2fdc4fd93ff660204;
mem[613] = 144'hff2efec300e5fe9f002201c3ff78fef4fe5c;
mem[614] = 144'hff84fe830092018efeacfceefe410314006d;
mem[615] = 144'h0153fc7bff3ffea40068fc7dfe16014f03e9;
mem[616] = 144'h00ef01900150ffaafeb7ffa2fd790057ffcb;
mem[617] = 144'h00fbff0f01f8fe29fda7ff6a00a6027c00fb;
mem[618] = 144'h041504270577fdfcffef01b2032e02de030b;
mem[619] = 144'h01de01f700a7fb020319ff9c066f01de06e5;
mem[620] = 144'hffbf0345fee8fc57ffc0ff24fee9033cfe68;
mem[621] = 144'h0211fe9801ee0b940db503a2fb7ef99b0194;
mem[622] = 144'h00b0ffb80126ffe40076fe2e00de00fc0013;
mem[623] = 144'hfddcfe9f0033004a00f6fdc2fe7bffb00166;
mem[624] = 144'hfec4ff27fde70176ffe5ff89fed7005cfec4;
mem[625] = 144'hfeacfed3ff31fdfcfe4d00c7fdb3fe2200cb;
mem[626] = 144'hffe400a4feeffff9ff1d0044006e0101006a;
mem[627] = 144'hfe8cffe1fe5a0007009aff150129ffb50112;
mem[628] = 144'h001f00e2fdcdff91008bffd4fef9fec500cc;
mem[629] = 144'h0181fefd0167fe85fe4a00d8fff7fedffff7;
mem[630] = 144'h013bff5f007600fefe8500ca009e00070131;
mem[631] = 144'hffd0006e012efefcfe42fe9d003d0142ff0a;
mem[632] = 144'h0228fddbff9d0104004f00a5fe46ffee0198;
mem[633] = 144'hfe83ffc10129fe8000320013006d00dfff11;
mem[634] = 144'hff7efe93010000c201fa00cefeb7ffb1fddc;
mem[635] = 144'hffc1fe8c01100018fff100f0fdc000850025;
mem[636] = 144'hfeb9feb9ff08ff88ffee00a3fde7ff2100ca;
mem[637] = 144'h00d9019001c9fe970099ff84fd5eff88ff81;
mem[638] = 144'hfecb016f016e012000ee00ba0058fe7cff3d;
mem[639] = 144'hff61fec8ff8aff34ffea001e00b6ff1fff41;
mem[640] = 144'h0471038d063303bbfd68fa9f04eb023d02e7;
mem[641] = 144'h046f02f703abff7efea2fddb014ffd71fab1;
mem[642] = 144'h0014ffc3ffdf007cffc4012fffa4fda2f7bd;
mem[643] = 144'h03a904b903d6fc63faa2006d000d002affa1;
mem[644] = 144'h01e2020d046f0247001cfc5d04a802bf017a;
mem[645] = 144'h004aff2a008cff44fef2012201f0020affea;
mem[646] = 144'h043f030f05a0019bfe37fe5003d2ff0cfcf4;
mem[647] = 144'hfed9007d036f00f8fed4fd230743026aff47;
mem[648] = 144'h04c40279028a0053ff6afe0000edfd47fe2e;
mem[649] = 144'h05e50294059801f1019dfe1102a3fda1fd7c;
mem[650] = 144'h0023fb29fd1b052f0152ff87fc6efa18f233;
mem[651] = 144'hff6bfc92fe80047bfce5fe06fdd5fee2f9bc;
mem[652] = 144'h017a031000ccfa92ff3a012ffcb9f95bfab7;
mem[653] = 144'hffb803750b2c030afaacfbb3064710c30984;
mem[654] = 144'h053502cb05170022ff75fe2302cafc9ffce6;
mem[655] = 144'h024102c804d3037c0090ff6a0368ff7efdc0;
mem[656] = 144'hfffe00660091fed6fe52fdb500c601b400b3;
mem[657] = 144'hffb10038ff12feb20021007fff660142005e;
mem[658] = 144'h015701a0fef50128fe48fff30139ff5fffa8;
mem[659] = 144'h0000ff1401030205010a0149ff55005900c3;
mem[660] = 144'h020b019bffea00cc013cfee9ff83fdc9ffb0;
mem[661] = 144'h008a009e00c2012dffcdfe3500fb013601c5;
mem[662] = 144'h01b0ffa5fe9dff340162007effcf0053ff2a;
mem[663] = 144'hfe59ff2100d5fead009700aeff1f01b5fe7a;
mem[664] = 144'hff3d004000b4fdaeffffff85fef0003800a1;
mem[665] = 144'hff10ff5500f6fed6ff4a004100edfe38ff41;
mem[666] = 144'hfdfe008f00d3ff31fddbffc1fea0fed2010b;
mem[667] = 144'hfdd7005701e7012a0126021aff93004b0269;
mem[668] = 144'hfe12016e007dff24fe570014fef60073000c;
mem[669] = 144'hfe1300a3fde6ff28fef9fffc0027ffa900a6;
mem[670] = 144'hfee5ffc300a8020a00fd00c800f300bafe67;
mem[671] = 144'hfe2a009f009cfdb1006c00950115fdf4ffa1;
mem[672] = 144'h01f5ff26fe1ffebcffe9fd2a052800bc0232;
mem[673] = 144'h02a601b4fef200440081fecf0071fdd7ffc5;
mem[674] = 144'h00ff01350183029700260124ff81ffb60102;
mem[675] = 144'h004bff1ffdedfcf8fe86ff4f0098fe8a00b5;
mem[676] = 144'h02bb035600f1ff1c0016fb8504530368035f;
mem[677] = 144'h018eff5100570076009702270058fed00202;
mem[678] = 144'h05bf008d0286fe9affc6ff31043bffedfe41;
mem[679] = 144'h0070fea0fc68fd10fdfffee2025602bb01a3;
mem[680] = 144'h036f02e0001501c000edfda6ffd000a601f3;
mem[681] = 144'h05e40368ffc40024018cfcb60113ffcc039f;
mem[682] = 144'h00cfff9503a801d3029a0275ffcff9eef281;
mem[683] = 144'hffeefe69fc03fe380003fff100b3fa3cfb42;
mem[684] = 144'h00bd008dfdf4fdc600270273fd2ffd46fee1;
mem[685] = 144'hffa001d005a60000fab0fdbd060c09be05b6;
mem[686] = 144'h02df0017ffb5fddbff36fe1202d4ff81fdae;
mem[687] = 144'h01800177013bff4dff18feef012900600292;
mem[688] = 144'h004a00ec02a30216ffd3fdb4ff70ff6200f5;
mem[689] = 144'hff2ffde100950086fd09fe7bff5e00500087;
mem[690] = 144'hfebaff4b00f00280013ffdc4016e039eff92;
mem[691] = 144'h030901ff0094004bfe38fc92ffd7ffa00043;
mem[692] = 144'hff09fec8011101e80199ff37001ffefaff93;
mem[693] = 144'hfdceff4afc55fd71fd7bfdf3ffa9fe11fd1b;
mem[694] = 144'hfefcff3aff8102d7ffd3fe23ff5dfebd00e8;
mem[695] = 144'hfff100f8fd5401a6ff7eff080255034ffeca;
mem[696] = 144'hfe97ff08ff87fef7ff69f9a6021fff54fefe;
mem[697] = 144'hfe970000ff070077ff32fdc2ff59fece0054;
mem[698] = 144'h0099fea1fd560609024403a4007efd22f531;
mem[699] = 144'h01aa0042feca04bd010e0416fefbff5efa83;
mem[700] = 144'h00affe9701c400a1faacff9702990114fd1a;
mem[701] = 144'h01c606f609fbffb103b2050c0203053702dd;
mem[702] = 144'h01dcfd78fe7e024bfcc6faab021f00240060;
mem[703] = 144'h0272fde3ff7700cdff7cfe65002afea900a0;
mem[704] = 144'h01d2feacfee202e401a301a8fea9ff940000;
mem[705] = 144'hffe3fd2dffdb0253feaffc9fff1d0123fd9d;
mem[706] = 144'hfdd8ffd4ff5fff77fe20fda2ffb7013ffd09;
mem[707] = 144'h0048fec6003a0489ff0aff44fe7f01780145;
mem[708] = 144'hfef4ff49fdc4ffcf028500bafd0aff12ffde;
mem[709] = 144'hfdf7fc23fc75fbe7ffd1fd21fe76fe24fcfe;
mem[710] = 144'h0172feca00bf026800b8fc97ff0d0084008c;
mem[711] = 144'hffc700ec00a702f80223fdb8006e0003013b;
mem[712] = 144'hfe1dfefe00e80174fe44fe7b014b009efbb3;
mem[713] = 144'h0034ff340050036100d0fe51ff88ff7efe0c;
mem[714] = 144'hff4ffd6dfa03fc85fed7ff48fca1fc44fc14;
mem[715] = 144'hffa4ffadfb63019f002ffe5bfe99fe720193;
mem[716] = 144'h0000fc56010502e1fb92fdf7019b01e0fca5;
mem[717] = 144'hfff9fe4dff93fc5601390009fd63fbac0050;
mem[718] = 144'h01a40130ffab0086fe79fbf9fe400108002a;
mem[719] = 144'hfe4bffd700d40222fe30fcedfd61ff8b0096;
mem[720] = 144'hfc90ff5401cfffd8fdb40200feb301a0fffd;
mem[721] = 144'hfe26001a00990050010f051c0101029702ec;
mem[722] = 144'hff7f02450284039b0444043d038900d9fd32;
mem[723] = 144'hffa1018e00e9fc3fff3a022a009501f20055;
mem[724] = 144'hff0f00d2ff6e021efe9b01db004101f502b9;
mem[725] = 144'hffcdff5dff1b007d00d6ff31001401a60299;
mem[726] = 144'hfcc1fdc002d1008401e103bcfe5b001b0174;
mem[727] = 144'h025efd4202cbfefcff820131fd53ff0b0171;
mem[728] = 144'hfc66ffef0315ffb8018d06d802ca04a10240;
mem[729] = 144'hfd87fdaf006600e10003026a002404560422;
mem[730] = 144'h026b02fefea2ff65012c01c000df0206054d;
mem[731] = 144'h012c00aafea6fe8bff34ffa202eb03af0594;
mem[732] = 144'hffc201520023fc80048101eb034402b900a3;
mem[733] = 144'h0063fee3fcc5047afe79ff12ffaafab8fd91;
mem[734] = 144'hff2cfdaf0283012c02af040000b6028301bf;
mem[735] = 144'hfe5400fd01c5010e0128041bfe88032602c6;
mem[736] = 144'hff95ff1ffeeffe0b017e0082ffb2fe9f0009;
mem[737] = 144'hff4201a400bfff730010fe9001830122ff5e;
mem[738] = 144'h010cfe7cff9f002affaafe5afef5ff61fe70;
mem[739] = 144'h00dc01c1ff38ffc201e0fee0001e013e009f;
mem[740] = 144'h00d5ff11fecffff5fed6fe6afe6300d400f9;
mem[741] = 144'hffd300b7ffeeffc900510168feaefe55017c;
mem[742] = 144'hff93009b013bfeef016a0005ff87fefefe46;
mem[743] = 144'hff71ff2aff620125012d0073ff5dff4bfe27;
mem[744] = 144'hfebcff2efeed006a0103fdd3ffd8fdcafffc;
mem[745] = 144'hfefafe82fde4013c00b7016cfe3ffeca0081;
mem[746] = 144'hfff0fdfcfebf01daffc20093010c018a0008;
mem[747] = 144'hfeae014a01b9ff1dfe8c0114008efefe004b;
mem[748] = 144'hff8dfddafdf70172fe4500a500c9fe38ff32;
mem[749] = 144'hfe57017cfe0b014800d9015dffcfff13fe38;
mem[750] = 144'h0185ff760194fec000a8fe980038ff92fe89;
mem[751] = 144'h002bff1d017700adff50012c00b0ff6a0176;
mem[752] = 144'h022f013403aa01f3ff160098030c00ff0142;
mem[753] = 144'h025c0235050afeb6017701ad00a1fe6eff44;
mem[754] = 144'hff6802c9ff42ff28008a026ffe300023fc86;
mem[755] = 144'h00bf01be029cfd6dfd080359014402dbfe49;
mem[756] = 144'hff8b012f03150409008aff710274034b00fd;
mem[757] = 144'hffbb0101019c00d90194fe6a01f5fea5002c;
mem[758] = 144'h00250207058aff490059037e0129ffecfd3c;
mem[759] = 144'h00d1ff4a02fa040bfe4e01f5036f025001cb;
mem[760] = 144'h0271060404a9fe2301ef054dfd76005100af;
mem[761] = 144'h00aa02be03beff01ff070257fef4010fffbd;
mem[762] = 144'hffbbfc1ffe33ffc80105fe9b0123fd72ff06;
mem[763] = 144'hffccfbc200c80242022eff62fee5fd5d0267;
mem[764] = 144'hff9204380067f9d900c2013cffa4ff37f97b;
mem[765] = 144'h00e6ff6806830ae1ff5ffe3d04540c57050a;
mem[766] = 144'h014d02b20544fe1e0065043fff110119ffee;
mem[767] = 144'hffb60118055f019101b30382010f02a2ffae;
mem[768] = 144'h024702c201b7ffe1ffb500ca02140184ff0f;
mem[769] = 144'h027802eeff21fe10010cff5c00cd0141feec;
mem[770] = 144'h016e0205004dfe02ff410159ff81014b02a4;
mem[771] = 144'hff8f035afe0e002500b1feb2039700abfe9b;
mem[772] = 144'h005803d001bcff9dfe54ff0f006c01170297;
mem[773] = 144'hfeda01e4fe6900bdfde6024a005ffe59ffff;
mem[774] = 144'h01be03d7026dfd000072ffbb01abffa5fd6b;
mem[775] = 144'h013f016f02870024ff2c014c02c001b40203;
mem[776] = 144'h02cc0346feecfe07ffd4fcd401700186ff3c;
mem[777] = 144'h020a042dffedfef500c200b702d7019b02be;
mem[778] = 144'h0069fdd8010b0210000002c8fd5efed80078;
mem[779] = 144'h0115ff9d023101310107ffea00d5034000f5;
mem[780] = 144'h010701e2fec6fff90210ff2cfedf006cfa6b;
mem[781] = 144'hffb700340590023bfd91ff780459070705a9;
mem[782] = 144'hff5a02240092fdf1fff8fe2f0231fffbff21;
mem[783] = 144'h004803b1014efdf8fea6ff370182034b01cb;
mem[784] = 144'h01f302b302bb02bf04610121fd16fcfffe5b;
mem[785] = 144'hfe59ff4cfee70199003ffe4dfeca020fffca;
mem[786] = 144'h0119fe72017efea2000100980050023a008a;
mem[787] = 144'h02ddffb00334053c02620023ff11ff5a0423;
mem[788] = 144'hfe8afff4fed2014801fc020e0163fd9afe9c;
mem[789] = 144'h002bfcf5fd7efdf3ffccfce1ff6dff8efef7;
mem[790] = 144'h0011fcbdff66005dfe08fefbfd730065fe9e;
mem[791] = 144'hff3d00db009903b3033700a1033900c2001c;
mem[792] = 144'hffd4ff3cfeecffe0feb5ff35ff83ffa7fe3a;
mem[793] = 144'hff5bfcf7010b01530152fe86fe5300e6fec0;
mem[794] = 144'hffd30056fc5d028a0154ffc801cb02d3ffb2;
mem[795] = 144'h000302bd02de03c701fa0250011001f0ffb8;
mem[796] = 144'hfeaa0028056200ddff3f0292014a02a001bf;
mem[797] = 144'h029e0465047800f006e905ac0027ff1dfde8;
mem[798] = 144'hff39fd98ffa802060071fe55fe4601eeff2c;
mem[799] = 144'hff45004b01d3014b02f9015ffe340062000f;
mem[800] = 144'hfef501beff1b009effd9fe0efda5fef3ffec;
mem[801] = 144'h0184fff40110fe17fd05fe34ffe7ff52ffed;
mem[802] = 144'hffabfeb0fef8fe90ffb2005000e300c20065;
mem[803] = 144'hfe1bff80fe3bfef6001cfec1fda2ff8fff16;
mem[804] = 144'hff64015100f1ffb2fe8bfe54fe9c00baff7a;
mem[805] = 144'h00acfeadfe5e019600e201a0ffcdff520132;
mem[806] = 144'h0036004afe6ffd52ffb80120fe7d011300b3;
mem[807] = 144'hfdc8005afe24ff71fd9800fafda8ff56fdd7;
mem[808] = 144'h002cfeb8fe8fffe6ff07ff79ff60ff140080;
mem[809] = 144'hffcafe69005dff89ff02fe96ff0fff9dfd77;
mem[810] = 144'hfed4fe81ff2bfead00a600d2ffd2017b00cd;
mem[811] = 144'hfd85fec1fcf60119fe79fe8efdfb001dfeef;
mem[812] = 144'hfe3ffe87ffef002dfe3bfff5ff8300980008;
mem[813] = 144'hfd86006601300083ffebfe6dfdcbfd47ff26;
mem[814] = 144'hfdc5ffcd0033fd74fefffe0fff23ff8bfe31;
mem[815] = 144'hff24012cfe4100c2fee6fda000b1ff1cff38;
mem[816] = 144'h0288020800c00133fe53fc70039702eaff27;
mem[817] = 144'h0214ffdefdc3fbebfde3ffbe04ebfd6bff7f;
mem[818] = 144'h0087001c0137fd2bfebeff050256ff9b0501;
mem[819] = 144'h01e3006b02bcffb3ffc0001d02eafe8b00b1;
mem[820] = 144'h041200ff00b9fd57fd25ff0606bd0449022a;
mem[821] = 144'hfebbff4d0059fd78ff74fddffea2ff110057;
mem[822] = 144'h038f034401300123ff63fbe90509ff0200af;
mem[823] = 144'h031e04b500e200c4fd70fdc40554036ffe73;
mem[824] = 144'h048c02ceff57fb72fbe0f9e80441fd2c0217;
mem[825] = 144'h059f00cb0164fe17fe9efc4c033d033fff8e;
mem[826] = 144'hffa2018509480818021303ccffe9010ef94a;
mem[827] = 144'h003103f804b9045cff33ffb5008a01eafaad;
mem[828] = 144'h0090009fff30fe3703d4017b0229fc72ffdb;
mem[829] = 144'h01ce046808e0059006bf03f4038209780453;
mem[830] = 144'h0460004c015cfd8dfd7bfdd4028e006ffdf9;
mem[831] = 144'h03b900e80134004afc41fbbd0631000efe7c;
mem[832] = 144'hfc9bfddcfef2ff17ff5903defd1b0099feb0;
mem[833] = 144'hff5bfb74ffed022302630217fff902660265;
mem[834] = 144'hfe17ffdd0291030b0106feba0077038afffb;
mem[835] = 144'h00ac0084fe1b02f40718ff6400d1011d037f;
mem[836] = 144'hfeabfeaffe6dfd16ffac0088fe1600daff24;
mem[837] = 144'hfea200070006ffaefeaffe06fee7032c0234;
mem[838] = 144'hfca2fe79feed01b50361002bfcedffd60314;
mem[839] = 144'h012f00e0ffa2ffac01c3004bfac7fdac016f;
mem[840] = 144'hfbbdfe12fe93002a01de003600e703be03ec;
mem[841] = 144'hfdb8fbdbfbedffcffe88ffe501e501650476;
mem[842] = 144'h034b01ff036000fa00560191014f05660629;
mem[843] = 144'h00e0061e014d018cfe2e004d01bb016200a7;
mem[844] = 144'h01a5fe3b04ea063303bfffb100ca04e5076f;
mem[845] = 144'h01e8fe77f67bfc5101bf02ecfc79f57bfa32;
mem[846] = 144'hfe25fd70fd0bff68031f00f4ff46008003bf;
mem[847] = 144'hfd47ff4efe34ffdaff6d000a009dffb10168;
mem[848] = 144'hfe2c018dfdbffdb903180305016102f1ff78;
mem[849] = 144'h00d301b5fb03fc2fff6f00a40010007b019c;
mem[850] = 144'h0168fecbffb6fcb5004700d9ff0ffdda090b;
mem[851] = 144'h010b023ffdce01a902d401dd01c90253fc75;
mem[852] = 144'h019502bfff7afd8cffe801a6ff9400da00eb;
mem[853] = 144'h00d502a6024d03080284015e02c304f503a7;
mem[854] = 144'hfed8031bfe39fd3bff07021b005202460120;
mem[855] = 144'h0173ff620292fcbf016cfff9fdfcff5d00c9;
mem[856] = 144'h023401c9fd46fce3fea901f902a6023903ef;
mem[857] = 144'hfec203c7fcd4fbfc00c30385021300ed0425;
mem[858] = 144'h00cc04ae0b3efe9dff12021c01bd06890a07;
mem[859] = 144'hffa103ae0793fa6d024cff3701b204c006a6;
mem[860] = 144'h009affbffce003340755009a031c02ce0259;
mem[861] = 144'hffd2fd6c01a30db10c3303b6fe54f8a1fb21;
mem[862] = 144'hffb70019fcfafe5afebb0290022f021c00d9;
mem[863] = 144'h0126012dfe55fd7601750303002502af0119;
mem[864] = 144'hfe970308018301970011fd44fe6cffc80163;
mem[865] = 144'hffe902e8000e01b8ff0cfdcafed9fe240182;
mem[866] = 144'h00f7ff11ff760145ffbd0170fddefd41ffe9;
mem[867] = 144'h005e026c020eff80fcf4ff020061fed403a0;
mem[868] = 144'h012a027900660260010bff49010dffe7ff85;
mem[869] = 144'h034f00130200038301bc041e034e003d015a;
mem[870] = 144'hff7d003f0009ffdcfe02fea5ff76ff42016b;
mem[871] = 144'hfe70ffa9fea1015e004bff0201b4fef60215;
mem[872] = 144'hfe6d001102bb0142fede007cfe27fd5800d8;
mem[873] = 144'hffa9ffff02380122019b00d2fc50fcc900c0;
mem[874] = 144'h0061002aff150276009201d003600114fed7;
mem[875] = 144'hffd7ffedff1900aeffaefffb00b8009cfff1;
mem[876] = 144'h0293023400d0ff910128fed9fd95ffb00316;
mem[877] = 144'h0196ff15ff5b00dafe03017603c402ce0404;
mem[878] = 144'hfe9302d302fa022b019a0155fcd3fefb01b4;
mem[879] = 144'hfe33002f024e0234ffe20070ff8b009eff83;
mem[880] = 144'h0132029f028001740323fe4afe3bffb60194;
mem[881] = 144'hfed902e50314ff6e0057feb7fcf4fe97feef;
mem[882] = 144'h00a7fff9ff87009002aeff54fc78fe4afc11;
mem[883] = 144'h010a01810175fff1fb13fd1d008500fffed9;
mem[884] = 144'hfe6700ef037203f201ccff86ffc6fe5f007a;
mem[885] = 144'h0098005e0033fe64ff4e01d30043ff66fdb9;
mem[886] = 144'hff7000e5029a008eff15ff33fd20ff3afeaa;
mem[887] = 144'hfd3600e903490218009dff3b0314ff0fffb7;
mem[888] = 144'h012c0381032703bc0180ffccfd42fcb8fccb;
mem[889] = 144'hfeb300aa04b104fd013801d4fbd5fd29fd51;
mem[890] = 144'hfd85fceffc5afd35fd9a0142fff9fda3f923;
mem[891] = 144'hfddcfc9afe6fffbc00930286fff5fe5ffd1f;
mem[892] = 144'h0189017300affd26fc43fdfafe99fecafad8;
mem[893] = 144'hfe8b0079043e0209fc0dfcb2032a0a1b0633;
mem[894] = 144'hffa002310355001800240038fde6fd3ffefc;
mem[895] = 144'hffae03d202e4041e03a8feaafd58fe79ff7b;
mem[896] = 144'hff96fcaefa84fc9efd3f013affe1fd66004b;
mem[897] = 144'hfdbffbeafddbfeac01320293ffd2feae06c9;
mem[898] = 144'h01a2ff56005e031a02db03c9003000fb0631;
mem[899] = 144'h0012fb26fc3700b901510098fd20fcd60420;
mem[900] = 144'h013cfdb8fac2fb5bfcee0042001afefafe9f;
mem[901] = 144'h030a020a026602fdffab0294ffef026b0338;
mem[902] = 144'hfee0fb4afd09ffe7fffa0124fdb8ffb00312;
mem[903] = 144'h01c1fcb2fb4efd57fe01fed8fd18fc8a0034;
mem[904] = 144'hfc67fc46fdf9fe7c018801f9ffe4ffae0496;
mem[905] = 144'hfec7f904fa52fd79fe9b008d00d7ffb90499;
mem[906] = 144'h03b008d80780ffa8ffed03d1053b0492f92c;
mem[907] = 144'h045c0489fdb3f90cfdddfec5034bff28fb62;
mem[908] = 144'hfe39fc2e0120ff60ff5d02c6007900e208b5;
mem[909] = 144'h03d3059102cd06c507dc03cf0144fb66fce6;
mem[910] = 144'hfe47f951fb2bff97ffe00362ffd2fe130455;
mem[911] = 144'h0009fd95fce0fe130194ffce004eff0a03a9;
mem[912] = 144'h009efed1fd9bfde1ff49fda6ff5700a9fe63;
mem[913] = 144'h00ff00b1ff6700a9fe6afe2dff74ffab00d1;
mem[914] = 144'hfe8cffd4ffcbfe4eff0a0054ff21ff9b007b;
mem[915] = 144'hfddbfd98ff56ffe1ff9d010bff0cff7e0116;
mem[916] = 144'hffc5fe04fe74ffcb00a90088fde5fe4dff1b;
mem[917] = 144'hff4a012efe89fedd016afff7002a01c0ff5c;
mem[918] = 144'hfe9b008ffe6eff35ffe9ff960023fe6c0036;
mem[919] = 144'h00df0074011900510090fffe00fdff73fef7;
mem[920] = 144'hfe7dff8afe3c0025fea4002cfdd80127feec;
mem[921] = 144'hfdeaff6dff7cffd9ff8eff04febdfdf1fe66;
mem[922] = 144'hfebd003dfeb300f300670050ffa2fea00102;
mem[923] = 144'hfef3fdf1fd98ff550078fd76ff12007cfe2b;
mem[924] = 144'hfdd2ffb7feacfe9f004ffe6efdceff2100e6;
mem[925] = 144'hffa9fdc8ff17010500fc0138fdae009ffe2b;
mem[926] = 144'h0093febffeea0101fefdfefafde400f4fefa;
mem[927] = 144'h003dfdf0ffab0009ff4fff6bfd8a00f700ff;
mem[928] = 144'hfc7efe05fe8efecf004301d8ff23043d016a;
mem[929] = 144'hfe85017100aa01e1014200f5ff8d03f402b0;
mem[930] = 144'hff9dff4502e80284007801c8ff770233fe9b;
mem[931] = 144'hfe0d01c4001cff8efecd00e001b90264ffe6;
mem[932] = 144'hffd6012a0120008d000301d4fd4c01540295;
mem[933] = 144'h017b00a4ff7efdf9fd95001500e300ac0152;
mem[934] = 144'hfd2302000122012500d3027bff7d036d0312;
mem[935] = 144'hffdffecf027afea1ff26ff69faec00490219;
mem[936] = 144'hffbb0299010801a20138035d0234056b020b;
mem[937] = 144'hffe80189006e0221ff620274012902f501e9;
mem[938] = 144'h007bff13fcebf9c8027fffeafc59fb5e02fa;
mem[939] = 144'hfe47fd46fa17fe04fe52ffd0fdcefe2806eb;
mem[940] = 144'h013d00170083ff59fe6aff9501c403e4fd8c;
mem[941] = 144'hff7bfdc5f946f8b4f772fc5dfd28f78bfe18;
mem[942] = 144'hfe200117017dff8b00ab019700fb033d04b4;
mem[943] = 144'hfdf1ffc4013b018fff3a02bcfe45048d012a;
mem[944] = 144'hffc200cafd65fe1ffdacfd890076fe9bfd77;
mem[945] = 144'hfe9d00e800adff8d0086fd68fe4afe84fe5e;
mem[946] = 144'hfdd7fdaefd86ff68ff14ff4cfe25feb2fe03;
mem[947] = 144'hff17fe0efe3afe6a00f5fe0d00bc0039ff69;
mem[948] = 144'hff8bfdefff58fffeff4afdc600a4fe69febd;
mem[949] = 144'h005d00dc002101cdfe1fff89019e00bbff36;
mem[950] = 144'hfdfefddcfe47fddffeb2fe51fda1ffe5fda9;
mem[951] = 144'h00be0123fdb3fea7fdebfddc001000be0026;
mem[952] = 144'hfe8dfe2affd0fe60ff00fdf8fe41fe7bfecb;
mem[953] = 144'hfeb6fe9dffaafdc8ff9ffdf10039fff1fedc;
mem[954] = 144'hfd7bfd7a00e3ffc2fe03ffeafdff006e00d3;
mem[955] = 144'h00c3012bfdbeff97fe3cfe33ffa5fe6ffd5e;
mem[956] = 144'hfdb0ff20fff2ff58ffc5feacfec6fed4fffe;
mem[957] = 144'hfe47006bfdb0ff8dfe77ff7cfe50fdabff01;
mem[958] = 144'h007ffe70ff05fe28ff0aff0a00d2ffba005e;
mem[959] = 144'hfec8fe7afde6fe940091ffd4ff75fe170063;
mem[960] = 144'hffec0114fe48003a001fff54fe56005aff1a;
mem[961] = 144'h00c000eb00f4fe73ff06004ffe9ffff8ff73;
mem[962] = 144'h018e01080047fe7000e6fee900b8002fff82;
mem[963] = 144'h0100feb6009400d1ff9afe7cfff20148fe59;
mem[964] = 144'hfed40025ff070037ff5b00e3fde4ff4afef8;
mem[965] = 144'h00c8ff5e00700189ff52fe27ff22ff2eff0d;
mem[966] = 144'hfe2bffb000af0150ff25fefdff40ff23fff0;
mem[967] = 144'h00a7fe80fe8e009bfe73ffd9ffaefec401bc;
mem[968] = 144'hfe61fe6ffdbdfe0afeb8fe690096ff6dffa7;
mem[969] = 144'hffbaff23ff86ff82ff210030ffc4fdc7fef8;
mem[970] = 144'h00160148ffc7006eff4a0171ff07ff8efe86;
mem[971] = 144'hfdd601670094ff88ffaa00dc0037feebff02;
mem[972] = 144'hfef8ff020098fddefe60fe6200ab00edff28;
mem[973] = 144'h013afe960129fde400760093ffd300beff99;
mem[974] = 144'h00d3005c01b0000b00b9fe5b0026fe3dfee9;
mem[975] = 144'h0093ff8f007600c1fe7bfff8003c0177ff62;
mem[976] = 144'h010dfd0d0200fe99fd1afd1fffa8fe25ffac;
mem[977] = 144'hfe29ff52fd50fdedff65fce0fd66fde1feb2;
mem[978] = 144'h008efe2b003bfd99fcd4fd1400380079fd3a;
mem[979] = 144'h01eafe7002ebfcb0fe9eff0f021cfe38ffd2;
mem[980] = 144'h008a015202520004fd5efdc3022901ccff3f;
mem[981] = 144'hff99ffecfee10015ffd6002b003dfe24019a;
mem[982] = 144'h0011fccb0080001bfeca00060188fe83fd33;
mem[983] = 144'h008100c7025c02ac0004fe2effb2ff77ffac;
mem[984] = 144'h020eff5ffe0cfdf7fd900001ff04ff82fd3f;
mem[985] = 144'h0004fd0dfd39ffaeffc2fde90223fe7ffee2;
mem[986] = 144'hfd65fd960060024effb5fd4b0067fdcd033a;
mem[987] = 144'hff5dfe22002c02dbfdabfd08fd06ff8f00f7;
mem[988] = 144'hffd00034ff9ffd8300a0fdc9fce7fe73ff3a;
mem[989] = 144'hfd1c0002fe58fee6ff54fdcbff04000c00a6;
mem[990] = 144'hfef5fd430032ff38fca1ff10011cfffefde2;
mem[991] = 144'hffc1ff55fe9e0061fd16fe270232fe36fd8e;
mem[992] = 144'h03ae015002c40210028c02f60061fcc9fec4;
mem[993] = 144'h02da01a3fe8ffdcbffa8fdf8fdc2fdc2fdd0;
mem[994] = 144'h0024fcd4ff59fd81fc5bff09fef30080ff35;
mem[995] = 144'h0240002b00ba04bd030f01ecff6fffeafe07;
mem[996] = 144'h005802020235001d03c1015202bd00aaff83;
mem[997] = 144'hff95fde3ffccff93fc93ff2afd26fef6ff9c;
mem[998] = 144'h0353000efdaefd11ff3bffe0015ffd72fd80;
mem[999] = 144'h01cd04dd017401220377016a0628028dff61;
mem[1000] = 144'h03df002efe42fcbeff3ffd24fdaffcaffdb7;
mem[1001] = 144'h04470035fec6ffd8fe61fe23fe37fc1bfce0;
mem[1002] = 144'h0065fdd1ff08051701a1feaa00c500ef00e2;
mem[1003] = 144'h00e901a905eb055c012b022c01f903870098;
mem[1004] = 144'hffe5ff4601d004a603ad032cfddbfe5602c1;
mem[1005] = 144'h00a1038207120059029b04ac038f06befeb6;
mem[1006] = 144'h046300f8001f00f5fe1bfd7c001efec3fbd6;
mem[1007] = 144'h038dffbdffb800a8fe12fdb70020fc97fc8e;
mem[1008] = 144'hfd8bfcb2ffd4fe37027001b1fdef010d04dc;
mem[1009] = 144'h00c80159017901ce031a035a010d02f20344;
mem[1010] = 144'h022f023c057f05c4028e0029ff8e00da0259;
mem[1011] = 144'hff21ff67fde0ffd1ffd70050fea002960036;
mem[1012] = 144'h0138007001b501a4019202b9feeafe870134;
mem[1013] = 144'hfea0fdfeffddff190018febf001a01140187;
mem[1014] = 144'hfd600165ffca00b1023400defdb200c00119;
mem[1015] = 144'hff04fd12fcaafe070086016bfbea00d7051d;
mem[1016] = 144'hfe79032602ba025102260307fe6f002f02de;
mem[1017] = 144'hffe5008e00d2024402fa0000fdbc0265018a;
mem[1018] = 144'h035d01fa0093fe8600a300f201fc006dfda5;
mem[1019] = 144'h02220045fd71f8b9fe9a01170223fd6703af;
mem[1020] = 144'hff5402d50169fdabff3000b900a2029d00d2;
mem[1021] = 144'h0178003dfbc7052d05240393000ffc710874;
mem[1022] = 144'hfeeefeb900290315002102e3fcee01c00286;
mem[1023] = 144'hffcd007901ab020b037101e7fe6b017801b9;
end

always @ (posedge clk) begin
	q_a <= mem[addr_a];
end

always @ (posedge clk) begin
	q_b <= mem[addr_b];
end

endmodule