module convolution(


);

endmodule