`timescale 1ns/1ns

module wt_fc1_mem2 #(parameter ADDR_WIDTH = 11, DATA_WIDTH = 144, DEPTH = 1024) (
input wire clk,
input wire [ADDR_WIDTH-1:0] addr_a, 
input wire [ADDR_WIDTH-1:0] addr_b, 
output reg [DATA_WIDTH-1:0] q_a,
output reg [DATA_WIDTH-1:0] q_b
);

reg [DATA_WIDTH-1:0] mem [0:DEPTH-1];

initial begin
mem[0] = 144'h0398069803a30176ff4d016d021903df047e;
mem[1] = 144'h02f305ac0497029affbcff79024a03b9017b;
mem[2] = 144'h01c704bc022ffeb701dc063e037a0116faea;
mem[3] = 144'h01ac01d1038f0331015600e60329014f010f;
mem[4] = 144'hffb7037803a70321006b015f01d000e5020a;
mem[5] = 144'h0038005f0097fcc4ffaefecb024e008a0058;
mem[6] = 144'hfe000235014bfedc00cdfddefe5dfc8dfc61;
mem[7] = 144'hffe4fe5f00e4ff8203670272ff3ef9cdf964;
mem[8] = 144'h030405a104320000000cff75005f018c0098;
mem[9] = 144'hff190373005600cdfc98fdfe001000e40235;
mem[10] = 144'h0204048405580235fe860024000402dc02a8;
mem[11] = 144'hff8a0326fca5fb11fc73ff79ffda06f6fb21;
mem[12] = 144'hfdb4ff97ff54ffecfde90150ff5affe40132;
mem[13] = 144'h01f10000ffb8015e01ddfe5effef010fff33;
mem[14] = 144'hfdf7fff5009702c4024301f8004902830193;
mem[15] = 144'h013a031701a0031a02710191007c03ee03f4;
mem[16] = 144'hfff2fe22fe2f00b2ff4fff30ff9dff5bfe91;
mem[17] = 144'h0095fec4fe9cfe18fe7c017500af0154ffcd;
mem[18] = 144'h00800217ff9d002d00a300bf007c00a8feac;
mem[19] = 144'hff68ffd1fe87ff7dfe73ff47fee0fec6fef1;
mem[20] = 144'h00170055fe4ffff9005f0090fe73fe27ff8a;
mem[21] = 144'h0010fe90014d00340061010d006aff37ffb9;
mem[22] = 144'hfe87021efef9ff970133017d0067006d00fd;
mem[23] = 144'h004101ae0179febe01360015fdf6fdf0fdbe;
mem[24] = 144'hfe16fff9fea2fe44ff3bfec6ff2dfe55fef7;
mem[25] = 144'h0191005dff8f0209fdc8ffa6000b001600f7;
mem[26] = 144'h0091ff83fe10ff7e00e90023ff61ff8f00b2;
mem[27] = 144'hfe030180022502110234fed7ffcafffe01e7;
mem[28] = 144'hfeddfe65ffd9004701c9006e00b3ff61ff8d;
mem[29] = 144'h01280153008601b40137feb3ff0cfec1002d;
mem[30] = 144'h00fc00fdfe320067004600d7ff75fe47fe2e;
mem[31] = 144'h00c4006e0095ff90fdef000300dc016bff0a;
mem[32] = 144'h003eff99012000840154000b0076fe350179;
mem[33] = 144'hff3f016e00d3ff23fe3700bcfebe00d40161;
mem[34] = 144'hfe81ff80ff20006b017b009fff3efe76007d;
mem[35] = 144'hff9b015aff04fe9100b600f7ff6afedbfffe;
mem[36] = 144'h017a005a0036ff780065ff0a00dd0159ff40;
mem[37] = 144'hfff0feb4ff120158ff8bffaaff27fe8bff9f;
mem[38] = 144'h0183fe5f017cfea0fdf4ff2afffc005aff39;
mem[39] = 144'h00fd0019000fff9dff560021ffbdffbe0102;
mem[40] = 144'hfed7fec20017fe19fe3dff95fde7fdeaffda;
mem[41] = 144'hfff7ff4e01ceffb9ffca0154fffbfff8ffb0;
mem[42] = 144'hfe86006afe3bfe46ff28016efefe01a90157;
mem[43] = 144'h0085fea2fefe017a0002004b00f900fb0199;
mem[44] = 144'h0011fe2fffc1018dfe3c0179010e0101ffed;
mem[45] = 144'hff9ffe46fe46012900ebff35ff5afe6dff03;
mem[46] = 144'h0085003f001efe53004dff7500c8fe820032;
mem[47] = 144'h005afe31ffe3fe7ffde8003a00a6fe5bfe87;
mem[48] = 144'hfdb2004ffdf300f6fdafffe0ff7200530019;
mem[49] = 144'hffa9fda9ff38febdff7aff4affa20081fe54;
mem[50] = 144'hfd8300ebffa700daff69fe3effb5fe13ffb3;
mem[51] = 144'hfe330085fec1fe8ffff7fddffd75feb9ff7f;
mem[52] = 144'hfd5e00faff74fe4cfd88fe88ffc4fe0bfdde;
mem[53] = 144'h008000d9fe0cff17feb1008700bffe5cffe7;
mem[54] = 144'hfd9cff4ffe78fd7800880019fef7fde90029;
mem[55] = 144'h01100053ff38fe58ff4300defe540058ff88;
mem[56] = 144'h006bfe65fda8fe8c003a00e7fe5affb9fef6;
mem[57] = 144'h00c40082fd6800a0ffbcff23fdb1ff9cfecf;
mem[58] = 144'h001c00bcfdf70066ffe2ff67ff45fd570024;
mem[59] = 144'hfdfe01a5ff8efecfff490018fdeefec6001c;
mem[60] = 144'h00f5fe79ff9fffc500f6fe32fe77ff970171;
mem[61] = 144'hfe8001b8ff12fe3f0138006afe76fe40fe80;
mem[62] = 144'h00c7ff83fe7efe34fe58ffc1ffe20053ffb5;
mem[63] = 144'hffcafe6300e3fde1fdc9ff8cfda5007bfddd;
mem[64] = 144'h04e803f302f7000300d0ff7bfd6f012ffd5d;
mem[65] = 144'h0346054c00ebfe1f0074ff62fe96fed1ff2d;
mem[66] = 144'h0503ff5ffcb5029900420147fee3fd6c0014;
mem[67] = 144'h04060208ff97000effa6febbfe02ffcefbd1;
mem[68] = 144'h03900557febf024cff43ff4efcec00affbc7;
mem[69] = 144'hfb89fdad0478ff3401c9fe230069042e04d2;
mem[70] = 144'h013cff41008c01eafc1cfe7dfc88fd50fd7a;
mem[71] = 144'h011bfb74f94d029cfa96fe0cfe43fbe8ff03;
mem[72] = 144'h044101f40101fec50004000dfe7cff59fd81;
mem[73] = 144'hff7b02490096ff0dfe23007afb56ffa6fced;
mem[74] = 144'h037d041b00a4003e0047fd38fb68fbf3fdca;
mem[75] = 144'h042afd01fce9073802eefd1701e8fe0703fd;
mem[76] = 144'hfe290100fef40087ff3dfe510005fd3fff3d;
mem[77] = 144'h0141ff33fe6dff0f0145ff9cffd80147014f;
mem[78] = 144'h00d5020f0256ff9e032501defea203a0fed6;
mem[79] = 144'h017904e1fe1bfee7fdeefe78fec7ff4eff82;
mem[80] = 144'h001cff28019700a20112fee7fecbff7fffe5;
mem[81] = 144'h004effb6ff40006300fa0135fe2800a8022e;
mem[82] = 144'hfe44ff680095fe2c00ee0024fddeff6f00f4;
mem[83] = 144'hffde01550138012900dcffbdff4dfe67ff52;
mem[84] = 144'hfee7fef700c8fe97fea3ff380180fe12fe2c;
mem[85] = 144'hff70fdd1ff6c010c0107ff0cfe59ff41fe42;
mem[86] = 144'hfe4e0168020101200130fec5ff9600790077;
mem[87] = 144'h016bfeca00dbfed3fe9cfdfcfecbfef30112;
mem[88] = 144'hff63feeafebaff8cfdeeff72ff8d00ef00ac;
mem[89] = 144'hff7fffe201070177008e0065017dff7800c1;
mem[90] = 144'h005f01d1feeafe7e009600f501ddff23fed2;
mem[91] = 144'h004efe94ff76febb009800f5015bff9600e9;
mem[92] = 144'hff80019afe6ffe7e007d0090fef8ff7bff48;
mem[93] = 144'hffd2fe1f00dafeaafec7feb7ff12fead01be;
mem[94] = 144'h0026ffe400c0ffc2006eff7afe75ff9c0084;
mem[95] = 144'hfe7afe53ff9dfed2ff09fedb0148fe84fe1f;
mem[96] = 144'h047103e10374fd77ff200334059003b303ea;
mem[97] = 144'h012504de045ffd4efd6b01d5059205a304dc;
mem[98] = 144'h045d061eff3bfe3c026e08d502830237fdd4;
mem[99] = 144'hfffe023d043afe0a00d50256026302b501c6;
mem[100] = 144'h00790421030c00f0ffd6017103d0021204b1;
mem[101] = 144'hfe46fb95074404c8ffaaffe4fddcff0d04b2;
mem[102] = 144'h02c602fdffe1007702da030102eb024e0284;
mem[103] = 144'h02b4063cff0ffeb2044c010b0234fbc6fb04;
mem[104] = 144'h02be01b601acfe90feb503c3039405a70475;
mem[105] = 144'h02bb00e1025f00b0fd08009a014c04a703b4;
mem[106] = 144'h03440370064a022300a60339033304e403c0;
mem[107] = 144'h051c00fdfe83fd4c03f0ffb0060d0559fe65;
mem[108] = 144'h02a1035001d100ccfeea003a02b6028d00a3;
mem[109] = 144'hff73fee9fe32ff1cfe57ff4c017ffe5c0058;
mem[110] = 144'h0052ffa70232fb68fdfb0360044606390630;
mem[111] = 144'h01fd037c04f6fd1900c401fa031b05eb0698;
mem[112] = 144'h000cfdfefdfdfe91fe8200eefef0ff3cffaa;
mem[113] = 144'h004e0047feb3017300c3fe6000760108ffac;
mem[114] = 144'h007f01ae016d00b2014cfed2009effe9000c;
mem[115] = 144'hfdcf0109fe290101fdff00fb013000e0fe7d;
mem[116] = 144'h0004febdfe7d00d5fefefe8afdec011ffead;
mem[117] = 144'hff420141ff64ff56ffc200cbffe6feeb0100;
mem[118] = 144'hfe350176ffbe01850099015dff96fe9d0046;
mem[119] = 144'hff6201560112ff00fefe015500d500c8ff88;
mem[120] = 144'h000b009dff520029ffc3ff5c00e0fe80fe84;
mem[121] = 144'hff390186fdf0ffa9ffbc00d70028ffe10168;
mem[122] = 144'h0125fe6800e5fef400600002003dffcf0155;
mem[123] = 144'h0170fec1fffa011dff37fe64ffe1016ffde7;
mem[124] = 144'hfe27fe8cff84ff9d01a7ff01009a016bfef3;
mem[125] = 144'hffb100ed01e200960053fe5100e00084ff7a;
mem[126] = 144'hfff1fddefffc001cfe76fdd30018ff42fdc6;
mem[127] = 144'h0059ff3700c1fe6800bdfea9fde3ff53ffe8;
mem[128] = 144'hfd56ffcf004e021702a7ff2afd30fccbffa5;
mem[129] = 144'hfd1eff84ffc102af0298fe76fca5fd72fd50;
mem[130] = 144'hfce6ffae00310346fb8ff6b5fc4d0082fd54;
mem[131] = 144'hfdfeff00fe09032600800199fcd30056006c;
mem[132] = 144'h014bfd16fdd1023e0351016b00040021fce4;
mem[133] = 144'h011e02ec0270fa9affce024f01bdffc403b5;
mem[134] = 144'h007dffae001400ca043f00b1ff2000c4ff8f;
mem[135] = 144'hfecf019201a9006bfafafa98024a0194fc9a;
mem[136] = 144'h00f6fcfbfef902720280ff26fbc3ff26ff3c;
mem[137] = 144'hffecfce6005e00ba01edfe45fe38fe8efd8a;
mem[138] = 144'hfdbffeccfd6dff10021f0036ff3fff29ff25;
mem[139] = 144'hfede01ec006a007fff4dfd04000f00da0377;
mem[140] = 144'h01d5fed5ff61ff6302030038ffc9fee1fed8;
mem[141] = 144'h010100faff0a019600760199011dfe5301a7;
mem[142] = 144'h03dc02ddff3d01c10238fef4ffafffae003f;
mem[143] = 144'hfe7ffe10fed1006701780084fb74ffc3fd40;
mem[144] = 144'h02eafcdafedeffe8010fff4a0662ffd1feb2;
mem[145] = 144'h03a1fe5cfcdbfe5802720178060700fcfd9f;
mem[146] = 144'hffcfff5ffd3800f703f303750120010d001f;
mem[147] = 144'h010cfd94ffb0feee020afff90432fe60005b;
mem[148] = 144'h0474fe70fcd4fdca0336017103830246ff06;
mem[149] = 144'h02130184ff86fd5801ee01cf01e9febff782;
mem[150] = 144'h03a1fcf0fef300f205b003f601ca02b00479;
mem[151] = 144'h02180117ff98066503a40658fe9802ad0462;
mem[152] = 144'h0247ff8aff12fe810256ff3e03ce0028fd48;
mem[153] = 144'h0421ff69fe8000e40480025d076d01dfffca;
mem[154] = 144'h03ffffb5ff3ffd9203ae0223062a004c00e4;
mem[155] = 144'hfc7d012afbba08320367fe73fd8cf9e4fc86;
mem[156] = 144'hfe92fd9bff3aff6eff01015301b600030039;
mem[157] = 144'hfebcffc10090ffda014a01c0ff86fe880104;
mem[158] = 144'hff9701cafe33fc30009a008d0526ff1efc34;
mem[159] = 144'h02e1fe50fc36ff56034f0254071c00c2fee3;
mem[160] = 144'h02b501150260005006a4023bfd2ffbabfd1a;
mem[161] = 144'h028d0377027ffe4f04c301b3fe68fbe0fe93;
mem[162] = 144'h0111fca1fcdd0a0bfe38fd0efd38fef5040b;
mem[163] = 144'h00620126fd6a015e0320ff24ffa0fd28ff8a;
mem[164] = 144'h00cd01e4fdea02dc04db005afe0efc68fff1;
mem[165] = 144'hff90fe5008e1fe5c028d01880234fc52f7e3;
mem[166] = 144'hfeb4ffad03030694fcd80127fd3dfece0419;
mem[167] = 144'h01f6fae903140ef8fa840040fe66015605f2;
mem[168] = 144'h002a04b3ff3f034005100067fddefc3dffc8;
mem[169] = 144'h0167026e00f2ffdf02eb0036fdf1fc23ffa2;
mem[170] = 144'hff2802520022ff440640ff83fc2efd54ff90;
mem[171] = 144'h0197fedaf9790e4601f403d300cdfc83fe1c;
mem[172] = 144'h002202afff7801d1fda7006aff4001680155;
mem[173] = 144'h0023ff9300c301b0016bffa4fe99ffe20181;
mem[174] = 144'h01210468018bff06052c011100cf004dfe76;
mem[175] = 144'h02290395ff2aff4a0300022d000afcb2fcd1;
mem[176] = 144'h00e1fdbeffd7fedeffe2fde6ff76febffea2;
mem[177] = 144'hfe9c0097fe53011bfedeff9601cf00ee0158;
mem[178] = 144'hff87010300db004500f0014afff6ffdf002d;
mem[179] = 144'hfe0fff20ffa2ffeafe560073ff43fe6f009d;
mem[180] = 144'h0070017bfef0ff52ffa4fdcaffbf00fffe9f;
mem[181] = 144'h014f0191ff5a0053ff4b015d00df011d01b9;
mem[182] = 144'hfdd1010fff1501b5fe6bfe780143fef3fe54;
mem[183] = 144'h001dffeafeb8ff3b0084012d00da0122fe90;
mem[184] = 144'h0123fec1fe56fea300a40173fdc000f7ff94;
mem[185] = 144'h01dc008101d7017a0033000f0205ff8eff4e;
mem[186] = 144'h0162014cff4d0094ff07fe0cff6101f6feb8;
mem[187] = 144'h00fdffbc012ffe8fffe9013e00ddfdf4ff0e;
mem[188] = 144'hff91014b0191ff1301680100012b00a3000a;
mem[189] = 144'h01deff16ff360135fe49fef300fbfeebfea0;
mem[190] = 144'hfed6fea1012affac017a012dffb1001400bd;
mem[191] = 144'h0018fef3ff58010b00a700aa00effeef000f;
mem[192] = 144'hffa7ff8601e0034701a5ff6afddb00f00021;
mem[193] = 144'h00f3015303410367fff1ff3d007f00ceff8a;
mem[194] = 144'h0382041f02ee0015fd1201890342017ffe22;
mem[195] = 144'hffab002402bf02b9023602290075013000d7;
mem[196] = 144'hfe470188004b03cd0131ffe4007ffeba0067;
mem[197] = 144'hfdd8f926fc7dfcb5fff5006c002a0695021f;
mem[198] = 144'h014404b8005f02f601c9ffcdfe85fd7cfdd3;
mem[199] = 144'hffd904bb0184fe04fdda00b3ffddfc77f83c;
mem[200] = 144'h0014ff1a030900f8ff5200be00cdff9f00e2;
mem[201] = 144'h0127fea800d2011300b0ff27fd58fcc3fcd9;
mem[202] = 144'h01b00270024202b202eafed2fdf4fe60fd78;
mem[203] = 144'hfff201ee01fbf789f5c2fc8201a402d00333;
mem[204] = 144'hffe5ffcefe14febf0225ffe4fe96000b00ec;
mem[205] = 144'hff22ff58fe6400e401ccff24ff94fe2bffdc;
mem[206] = 144'h00020136ff1d008202b30062fea9fe270041;
mem[207] = 144'h017e012c007601cb010b00dafeee006cff68;
mem[208] = 144'h0072ff7efe0602960070ffeffbabfb8bfaa0;
mem[209] = 144'h0138ff0800aa0334019ffe03f936fb0cf94b;
mem[210] = 144'hfcd4fa1602b706a1ff7cfe6afd90fb9f0269;
mem[211] = 144'h0069fe5d01d601c2fe26ff77fdbffae0fc82;
mem[212] = 144'h003dffb900a10425fefe0029febdfbe4fc9c;
mem[213] = 144'h0020046b001802b0ff6d011203d2014cff84;
mem[214] = 144'hfe1ffd15018e0035ff6400c70168fce1fd7d;
mem[215] = 144'hffd7fe6706030467fd76feaa0103020103e2;
mem[216] = 144'h007800c901060148029cfe41fc55facffc21;
mem[217] = 144'hffd4019bff7cfffb0219ff2dfb14fa0ef9eb;
mem[218] = 144'hfdffff31ff9a01bb023bffd6fc5ef9bbf869;
mem[219] = 144'h00cdfc4e01ae0a7304d7feeafef8fc7b0656;
mem[220] = 144'hff3100d9ffdf001fffb00083fee2015800b6;
mem[221] = 144'h002300ee00e5ff53000c01aa00d8fe57fe3b;
mem[222] = 144'h053203aafd9f040a0260fde6fc64fdb6fc94;
mem[223] = 144'h02070011fdd100fafeeaff00fa6ffa57fadd;
mem[224] = 144'h00850068fdf8fcdefefdfb75045f036cfe07;
mem[225] = 144'hfdd0ffa7ffddfe56fdb1fd59054b029f00a8;
mem[226] = 144'hfefb00380030ffb60063031d0321ffe5ffb0;
mem[227] = 144'hffb5ff73fe28fd1a0013fd0a01820067fedd;
mem[228] = 144'h009ffeefffa6ffd7007dfca4012a01ae001d;
mem[229] = 144'h01ecfdb9fd3b00440363fad5ff65fdf8faef;
mem[230] = 144'h007c025efff7fe3ffdeb01cb011b0260ff7b;
mem[231] = 144'h00ea000eff9901c9fe6f052cffdfff050031;
mem[232] = 144'hfe4eff9aff15fec0ffc8fc420529012ffe1d;
mem[233] = 144'h0117fe8affde0060ff0dfa0f052901e7ff92;
mem[234] = 144'h002701e8ff13fe0dfe9dfcd0035d03940115;
mem[235] = 144'hfb74ffbcf9ef0222fd910136ff69feccf9b8;
mem[236] = 144'hfd78005001b3ff23fe63fe430047fe76026f;
mem[237] = 144'h0136001400f6fe75ff1f01c10187fec301c6;
mem[238] = 144'hfcc1fc76ff28fefefef5fabb021b0016fcd1;
mem[239] = 144'hff270033ffe0fd7d017afb8302ea0170ff0a;
mem[240] = 144'h006103260217fc900090016ffec201530205;
mem[241] = 144'h03e6026902eefed6feba01a3fe4e0184049d;
mem[242] = 144'h00a7fe78f781ffd10231fc5afe85fe10007f;
mem[243] = 144'h012600a8fdf3fd9c00cc005f0158ff56023c;
mem[244] = 144'h016202b9ff9afe2402750245ff9c0106012b;
mem[245] = 144'h0384087d0d670011006d03ec0139ff82038e;
mem[246] = 144'h009ffed3fa09fffd0100f9f2fd14fe590586;
mem[247] = 144'hfe28fc1ff841049dff5af7270103fe7d0505;
mem[248] = 144'h016a01a0ff55ff1b01020052ff0b0318023c;
mem[249] = 144'hfc29020dff82fe2dfe50023afee3004a04f8;
mem[250] = 144'hfe60011801bbff4eff9f00d7fff8ff61024e;
mem[251] = 144'h04e601b5fefe074208ae074aff48023d000d;
mem[252] = 144'h019401b60090ff1bfdfbfffcfe99fe1afe0f;
mem[253] = 144'hfff0ffd7fe66019cff82ff5cfee6ff40ff06;
mem[254] = 144'h01cb02d3039dfbc3fdf90091fefe037f0183;
mem[255] = 144'h03b601b501f9fcdcffd902b6ff90ff940145;
mem[256] = 144'hfd37fd0cfece007a010200c5039202220257;
mem[257] = 144'hfca9fcabff7c020e0189000f04a000f501a6;
mem[258] = 144'hfd1eff85fc49f8e9fd9af7d703930055ff5a;
mem[259] = 144'hfe350044ff4eff21fef5ffd303c2036c03c8;
mem[260] = 144'hfe4bfc3600c3fd62021fffe6016e03410259;
mem[261] = 144'hffb5fc12f9c8fd2901d8040dfee7f85dfc93;
mem[262] = 144'h00e1fef1fe8effc005b6016d026a03ad03cd;
mem[263] = 144'h00120033fb4cfb1b0101fd9900e003050411;
mem[264] = 144'hfde8ffa101a2fec70149ffc502ae042203bb;
mem[265] = 144'hfe10fdc6ff5201c601620050081b0379033f;
mem[266] = 144'hfff0fd530003003c020201820377035c02ac;
mem[267] = 144'hfd6002f9fbcbf248fc8f015dfef6fe09f7e7;
mem[268] = 144'hff43005802d600ac027cff1d02deff9bfe53;
mem[269] = 144'h01660116febbffc000ddfe3c002a01af015e;
mem[270] = 144'hfdebfe0d02f600a7fc98fcae03690219019f;
mem[271] = 144'hfda4fdcf01bcff40004f0084031c022c029a;
mem[272] = 144'h03f502cb011ffd39ffce02f40026024e0491;
mem[273] = 144'hffdc03f903b5fc72ff5003be037804f0081b;
mem[274] = 144'h02280475ffd8018f0344047e011c0208ff79;
mem[275] = 144'h0266019a01f1fe82ffb6006a0195054b0200;
mem[276] = 144'h0108037a0322fe0d023b0240023c0247036d;
mem[277] = 144'h003700d409a501aaff8b01d4fe93fb51026c;
mem[278] = 144'h03290385025900bf0104fea8fe18011f028f;
mem[279] = 144'h030b024a01a502a10453fe56fec9fe57ffc5;
mem[280] = 144'h029a034c02d1fd1d017e02c101ee037606b6;
mem[281] = 144'hff360419040aff98ffc5033dfd6d053a05a8;
mem[282] = 144'h015903b4041efe3701430369ffdc03be0473;
mem[283] = 144'h027f027efd7102dc0788059302e0041bf883;
mem[284] = 144'h02a4ffac008c019cfda4ffcb01c8019eff1c;
mem[285] = 144'hff83000001baffbeffd6ff8b011bfe9e01cb;
mem[286] = 144'hfff10146ff1bfa3fff5903ef02af03cc062e;
mem[287] = 144'h004904a70284fc8affb803d2023d03220498;
mem[288] = 144'hfdd5fc95021203e80074fd7502690068fc7d;
mem[289] = 144'hfe5fffeeffb403e60229fdb50143febffb64;
mem[290] = 144'hff38fafffb84fb11fa4af88802e800bc013f;
mem[291] = 144'h0010ffd5016c005cfe00ff100354ff23fe74;
mem[292] = 144'h0088fcb200e501f3ffd8000f03e20097fc6f;
mem[293] = 144'hfecdf6cef583009604acffc5fc80faeafa46;
mem[294] = 144'h002efdf8fdccff67feec01ef02d10411ffcd;
mem[295] = 144'hfeebfd84f7cbf965fac4006d03d0028e04e5;
mem[296] = 144'hff9dfdd1019a0082fe2efe950364ff2bfbe0;
mem[297] = 144'hfef4fe4b004903650018fc4b030600c0fc31;
mem[298] = 144'h00bcfe59ff44ff7e0197fca004210231fc10;
mem[299] = 144'hfe50fca9fd30f660fbd10004ffd3f999fe78;
mem[300] = 144'h0230020100b3ff9601560103fe9100ac01a0;
mem[301] = 144'h0085fe5001beff4c0006004700fd0153016b;
mem[302] = 144'h004200c604c705390051fd0602dc0263fe3f;
mem[303] = 144'hfea5fee9015301c3ff6efba70069ff3cfd49;
mem[304] = 144'hfea7fed400140131ffa2fe3dff7afff2fe7c;
mem[305] = 144'h00edfecffe7ffff30146ff0dff9efe530084;
mem[306] = 144'hffd60108fd86ffc8ff31ffa40066fe810179;
mem[307] = 144'h00defdcefd94ffe800d90147fe92fec60122;
mem[308] = 144'hffe4fdf2ff73fe32ffe3fe0f007a00690094;
mem[309] = 144'hffa7fecffda2ff6dff27ffca012600e60148;
mem[310] = 144'h0096ff0dff79001efeff0092fe60ff900086;
mem[311] = 144'hfffafe4d00c6fdf8fe0c008b0009ff7cff8d;
mem[312] = 144'hfeb0ffb600c5fe67ff1c00950151ff31ff5f;
mem[313] = 144'hfec5fee1ffc3013a0050fe840007fe8eff69;
mem[314] = 144'hff35013efecefdd800b8feb4fe80ff62ff99;
mem[315] = 144'hff95fdd400abff0e002fff45fed6fe0cfdb8;
mem[316] = 144'h0130ff71fedffe9801c4ffcaff15fffeff7f;
mem[317] = 144'h00fb016bff2d008200b4ff90007b00f3fefb;
mem[318] = 144'hfe2800e400e6ff7cfdbfff2d0050fdda004b;
mem[319] = 144'h00220033ff57fefcfde9feb8005900670022;
mem[320] = 144'h01ea037102990087014f036cfb09fb550043;
mem[321] = 144'h03a60492027001d3042e02cffdcafccefee3;
mem[322] = 144'hfe95fdf0f8e80644043cfaddfb5bfbe30127;
mem[323] = 144'h026103c7fe7d010e02b0021bff72fbd4fdaf;
mem[324] = 144'h012701d200d001c40218020400e7fd0ffe08;
mem[325] = 144'h002107a209a7015b02a503a50500021afe6a;
mem[326] = 144'hfdf8fb65ff320194013dfca6fbdbfce50185;
mem[327] = 144'hfe10f713f9fc0554ff96f9e8fdccffd10443;
mem[328] = 144'h03bc033d0135018202d80126fce7ff2200bd;
mem[329] = 144'hfeda043c0206fe55ffb400bffbbafe80ff0a;
mem[330] = 144'h0074022afe720078034a00b1fc9efda3fd07;
mem[331] = 144'h03c1008f012f0a0f07050292ff2000d10420;
mem[332] = 144'h004bff5cff0c008fff8eff10fdf6fd5f00e5;
mem[333] = 144'h00dbffbcfef8ffe1fe8c0120ffc1000c0186;
mem[334] = 144'h02c7056b015e024002f903790040fe84fd07;
mem[335] = 144'h0056038300f0001f032bffd1ff0efe78fec7;
mem[336] = 144'hfd67fe7a0221009f04a701f1fc86fc72ffc6;
mem[337] = 144'h00ed00eb00660402040dff2cfc42ffc2fec4;
mem[338] = 144'hfe8efe4302840125fca2fa16fd99fffe0063;
mem[339] = 144'hff9efe9200aa044a022101abfe97ff0eff21;
mem[340] = 144'hfdcf00d10148046201430107ff14fefdfed0;
mem[341] = 144'hfe6cfd580028fa96023301e60034016eff9b;
mem[342] = 144'h017cfff8038601e3038a0229ff0fffcffcfc;
mem[343] = 144'hff4303650202ff39fc41f9ffffc20246fe68;
mem[344] = 144'hfec9ffd802bf00bb03f30104fdacfeb1ff1e;
mem[345] = 144'h00bcfe95ff800242027d0296fbf2fe88fe8c;
mem[346] = 144'hfed800260120043403430187fc74ff42fec3;
mem[347] = 144'h0122ffb2041ffd4afe06fe36004600630333;
mem[348] = 144'h002500fa00e2010e006e018b00e2ffceff45;
mem[349] = 144'hffd101280085012ffecafe890143fe430133;
mem[350] = 144'h038c0192020e034a01aa025cfe50ffb6006a;
mem[351] = 144'hfe8cfe2100fb0121037501e6fdd5fce6ff05;
mem[352] = 144'h0419019e0223ff01feca03c803ae0188fe4a;
mem[353] = 144'h02d00455013d019afea80311031a02fcffe4;
mem[354] = 144'h047501c2ffce02d40445069600ee0275febb;
mem[355] = 144'h02ba02270347046001ab050503240230ff95;
mem[356] = 144'h01a6014b025103b600ef046a007601670040;
mem[357] = 144'hfd84feb9040a0541fef5fe49ff8e02730142;
mem[358] = 144'h05e801ee030f044103fa0792feaaffa0fe5d;
mem[359] = 144'h046502c0ffd9063007e4068cff4affa0fd65;
mem[360] = 144'h02be01270369012d007a030203e502aeff30;
mem[361] = 144'h05c2005802f8ffdcfe0a0328ff3d00abfd1c;
mem[362] = 144'h032902f60236028f025c041b003effbc005f;
mem[363] = 144'h03a7ff83feb102d001da0042045bfc670209;
mem[364] = 144'hffa5fde600e801bcfdbdff8e035402d30150;
mem[365] = 144'hff78017eff9300aa012000effedbff7100cd;
mem[366] = 144'hff6b0186028a0024006cff7f0496027d01b6;
mem[367] = 144'h02bd0115007601110023031704c0025bff6e;
mem[368] = 144'h000fff8b000e01850029ffdeff0000befdc4;
mem[369] = 144'hffd3ff8ffe17ffa7015efe5cfdfbffd1feb5;
mem[370] = 144'hfe2b006afe69febdff210194015aff150120;
mem[371] = 144'hff47fef0fe14feab003afe7eff22ffd3ff4d;
mem[372] = 144'h00d2ff73013a00cf016afdd10167fe0ffe4e;
mem[373] = 144'h00fcfde9003b00a8001d017600370101ff1e;
mem[374] = 144'hffd9fe9dfecb0132fe250090fe01002100f9;
mem[375] = 144'hfef8007cfe88fe4afe2f0152ff9a0058fdef;
mem[376] = 144'hfe5a0169004bfe5fff7aff71013a0017fe0c;
mem[377] = 144'h015dfffe01d5007dff0bfec00054fe85012d;
mem[378] = 144'h01bf0158fecafe94fde60099016b0117002e;
mem[379] = 144'h005efeb9006a0014fe6aff8ffe05fe00005e;
mem[380] = 144'h01870020ffdcfe53ffe901710094ff400134;
mem[381] = 144'hfea9fe4d00b4ff0f0023fe23005dfed90017;
mem[382] = 144'hff56006c018100d5017e00b2fe30fdcdfe80;
mem[383] = 144'hff30014eff73fde1ff56ffdeffb6fed7fe64;
mem[384] = 144'h0231ff22fd5100a7ff090015fdd1fdccfd9d;
mem[385] = 144'h01d9fdfafcedfe40fe1efecffdcefdd8fff9;
mem[386] = 144'hfe5eff09fe42001d00cd00d4fe8bfdfaffc7;
mem[387] = 144'hffe9fdccfe48fdccff2b0000ff75fd03fe2a;
mem[388] = 144'hfe88fed2fec80026febc0110ffbbfd71feaf;
mem[389] = 144'hfdc202250043fddf0127fe1ffe6500ceff78;
mem[390] = 144'hff8dfdbcfe91fed5fea9fe5dfea2fd7dff57;
mem[391] = 144'hfd5cfff000b20168fe1bffbf0050fe92fef8;
mem[392] = 144'hff84ff14ff0aff0bfe07fd65fd8dfe70fcd2;
mem[393] = 144'h011800c9ffe1fe56002bfd47fcf8ff94fcc6;
mem[394] = 144'hfe67fff6fe18fdaf0039feeafd79fce7ffda;
mem[395] = 144'hff6a0020fdc0002402a1012afd8dfd61fe67;
mem[396] = 144'h00670181fe47006afeca007d011a0149fe38;
mem[397] = 144'h01ab00fa015ffeab009c01980174ff7301be;
mem[398] = 144'h0185feb1002afe89fe7e0022fe080086fe23;
mem[399] = 144'hffe8ff1efe9dffcf00cbfd16fe8efd8ffee9;
mem[400] = 144'h02e3ffe801b5026701ef00f00139fc86fd00;
mem[401] = 144'h0341034402870125035bfe480183ff40fe50;
mem[402] = 144'h03f0fc89fe9b059501b00618fe22fc5c0091;
mem[403] = 144'h032001a202190442010402930008ff8afe5e;
mem[404] = 144'h03d6014cfec603c5022effe201c6ff09fcb0;
mem[405] = 144'h009cffee024d01d80219ffd0017dfe7bfe2b;
mem[406] = 144'h0364016e02d804c3027c0648fe0bff7efd6d;
mem[407] = 144'h032dfec104c5060b025d03cdfe0801fd01d9;
mem[408] = 144'h043d0207016201900095025b00e5fd5ffe7a;
mem[409] = 144'h034702a301a2036f0089feccfe36fc52fd59;
mem[410] = 144'h049001a5fec1044f044d01b3ff11fefffcae;
mem[411] = 144'h03a2fcb0febc0a05fb6bff7c0083f9dd0472;
mem[412] = 144'hff76ff65ff5a00ebff2cfeb3010e01160102;
mem[413] = 144'hfe67fe21fff3ffd70117ffb0fe74005900eb;
mem[414] = 144'h020f026e019e02cc01e6fe560435039800d4;
mem[415] = 144'h01f60359ff9602d5010601d20142ff12fc55;
mem[416] = 144'hfe7dfd13fc62fceefc8bfd06fdedfdf3fd33;
mem[417] = 144'hfdf4fbeafcd7ff89fce9ff39fc0cff17fc4c;
mem[418] = 144'hff30ff3cfcd0fc52fe61fc78fc89fde4ff48;
mem[419] = 144'hfb95fee0fedefbc1fd4cfc7dfae7fef1fd4f;
mem[420] = 144'hfb79fc6bff32fea1ff70fcaefc51ff6d0068;
mem[421] = 144'hfe06fdc6fe71fe03fe0efdd0ff2cfb7fff99;
mem[422] = 144'hff05fe76fefdfc45fe2bff99fd5b010d00c8;
mem[423] = 144'hfd4cfe35fee6fbabff53fe0cfbe2feac02a0;
mem[424] = 144'hfe59fc16ff20fea8fed5ffb2fbd8fe5cfcdc;
mem[425] = 144'hfdf6ff21ff1bfebdfccc003afd3bff85fed9;
mem[426] = 144'hfe1efda1fc8afe2afd8fff21fa25ff050066;
mem[427] = 144'hfcf7fd90fff4fe33ff70fc54ff77fe64fc0d;
mem[428] = 144'hff8cff2dff79ff47015a00590130ff06fe99;
mem[429] = 144'hff4900ddffee00360160007cff83fe71fe48;
mem[430] = 144'hfcfefe53fe7b00d9fe4afd3efcaffd54fd8d;
mem[431] = 144'hfcd6ff42fd60fd96fd1ffc9cfc2ffd48ff19;
mem[432] = 144'hff55feef00b8ff36006dffcbfe310128006b;
mem[433] = 144'hfeb3fe1401b7ff27ff50fe1efe17fe48fe10;
mem[434] = 144'h015801de0072ffba0024fe6d009400210137;
mem[435] = 144'hfe5eff1aff79ff3ffea100b7008800a50159;
mem[436] = 144'h01570170011bff6dfe270122fec6fdf8ff61;
mem[437] = 144'hfde700a9fe14fe73ff17ffd3fea801080027;
mem[438] = 144'hfe79fee6fe1eff48ff53feb7fe6c003e0150;
mem[439] = 144'hfe75fda3ffc8fdd0ff39ffedfdcb00c7fe76;
mem[440] = 144'hfecfff8eff9900a000fd014bfeb1004afe35;
mem[441] = 144'hff8500ed003affd1ffb60119013ffe1f0006;
mem[442] = 144'h015efefe0177fe5000930131fe7ffe61ff24;
mem[443] = 144'hffa200380004fdac009a0160ffe2fec4fde6;
mem[444] = 144'hff04fff9fe41009fffce0055fe950116ff4b;
mem[445] = 144'h0032ff11ff7b01cbff9300caffddfe8e0063;
mem[446] = 144'hff94012fff9ffef5010aff7f00a1011c0152;
mem[447] = 144'hff97ffd0fe28fff4fe78010300adffb5fecb;
mem[448] = 144'h001dfffe0000fe5300eeff53ffd30023ff13;
mem[449] = 144'h0178ff2ffdedff42ff16fec8fece0105fdc0;
mem[450] = 144'hfece0094fdd8013ffe1900f3ff940025005e;
mem[451] = 144'hfe1d009ffe81014cffd3017bff5aff94ffd6;
mem[452] = 144'h0143013a0081fdfafe23ffac00f1ff07001f;
mem[453] = 144'hfee2ffd4fed7ff28ffe3fea0ff3ffeecfe9a;
mem[454] = 144'hfe03ffe40151fe18fed8ffb5011500bdff6c;
mem[455] = 144'hffff004bfe26ff2eff92fdc600d70068011c;
mem[456] = 144'hfee0fed90060fe35016affb000080083fe84;
mem[457] = 144'hfe83fe3a0009020301dffff4ffcbffa5ffb7;
mem[458] = 144'hffe900cffe3c0128ff91006500e7016f000f;
mem[459] = 144'hff4300a60006fdd9fe6d009e008800a6fea8;
mem[460] = 144'h0103ff11ff0301c5ff5f013ffe3600ae0181;
mem[461] = 144'h015e00cd01d8004d00b301a00141fec1ff3d;
mem[462] = 144'h00d000000062fff0003aff33fe82fde40046;
mem[463] = 144'hff63013efef90095001a0121004afe16005b;
mem[464] = 144'hfddb01af0206ffe60127011ffc7e0012024f;
mem[465] = 144'hfd8ffe2f01a60197ffa4fefffd5702e70368;
mem[466] = 144'hfd4a063c08c700fffa5207e8ff6a036fff8f;
mem[467] = 144'hfbd7020e02ac0477ff85ffccfdb5007a0271;
mem[468] = 144'hfdb9fedb052204a4ff59fdf5fe3b020c00f0;
mem[469] = 144'h01bbf9aafe5fff19fef3fd4300e3ff9b02ea;
mem[470] = 144'hfed106c0055f024cfc790008ff8afd26fc9b;
mem[471] = 144'h02200607076ffdbcff660433ff8dfefbf46b;
mem[472] = 144'hfacbfeef02f90340ff400177fcc900ca029a;
mem[473] = 144'h0025fd9b0225fee0ff5d0000fd84fd400246;
mem[474] = 144'hff080180046305370048ffa2fdcc001a01dd;
mem[475] = 144'hfb8303320432fcdff453fbe3fd95055a00de;
mem[476] = 144'hff2cfdd8febeff4d0156fe7400ae00af00ac;
mem[477] = 144'hff73febe0033febb005cfe2aff86ffbafe93;
mem[478] = 144'hfb75fe3bfe0f0027031e017dfbf4ffc802eb;
mem[479] = 144'hfcedfe44011a0215ff0b016bfc73016703e9;
mem[480] = 144'hf98f0219033501aafd5cfe11fa0201fc0369;
mem[481] = 144'hfbc9fc9f01500162fb88fd64fb0000a70208;
mem[482] = 144'hf9d20942089bfaecfdf407b4fe01046dfdd1;
mem[483] = 144'hfbe4000b05e9025ffc890110fd150111029d;
mem[484] = 144'hfe41fee40568038dfeef00ceff83025e002b;
mem[485] = 144'h01ecf8c8ffc70600fd1efe08058502310fa4;
mem[486] = 144'hff1906110596fbf0ff9502baff9efe93faee;
mem[487] = 144'hff5b05c105e2f7300593063d01b20124f567;
mem[488] = 144'hfa38ffd5062affe0fdc800e6fe1001f50310;
mem[489] = 144'hfc71ff05ff940080fbd6ffb1f940fc94fe50;
mem[490] = 144'hf96a005e050104d2fd17ff30fad0ff400044;
mem[491] = 144'hf9f004f003f4f658fc00fd01fd6609590773;
mem[492] = 144'h0087ffc90042ff76ffaafeabff2d0201fed4;
mem[493] = 144'hfe91ff3d01a2fe5b013efea6fe8afe5000e4;
mem[494] = 144'hfe0bfb52fe8e030effce0245fa45fef0034f;
mem[495] = 144'hfc94fd04053d01fdfd5affc7fdf20152042e;
mem[496] = 144'h01710114fe63fd990086fee500220002ff0d;
mem[497] = 144'hffa30022001effe4ff05feb500b400420043;
mem[498] = 144'h015c00dcfe110045ff44fdd2fec4fe1e0054;
mem[499] = 144'hfe0e0067ff9700c2ffa4fe86fe3000befecb;
mem[500] = 144'h00b4001c00aa005b0018fe99ff3e005bff10;
mem[501] = 144'hff85fe24feba0040012cfebf00b0fef1008e;
mem[502] = 144'h0018ffbffe58ff6900c6feef005b008dff90;
mem[503] = 144'h0046ffdcfdb3ff56fde6003c00c1fdc9fe6f;
mem[504] = 144'hfdd5ff35ff70fe1fff62ff7dfdce00dc0040;
mem[505] = 144'hff12ff770134feb2012b0006007b02270006;
mem[506] = 144'h00bd000300d501510118fdccfdfafecd0051;
mem[507] = 144'hfec9ff04feceffef000d01b6ff0f01a60044;
mem[508] = 144'hffa7018200d9fe9bfe2700a8ff9101dbff4e;
mem[509] = 144'hfeb9fe9d00ef0161016d00fdff7f01100106;
mem[510] = 144'hffcb007eff7efdf900c80072ff2900e2fee8;
mem[511] = 144'hfdf8fe35fdf2ff40fe530120ff80ff8afea3;
mem[512] = 144'hf96efd82fd920252fed9fe53f7d2fcef0323;
mem[513] = 144'hfb97fc79ff41024c0099fe1af931fbe20370;
mem[514] = 144'hf7d501540a87016efe260647fa1d02fcff49;
mem[515] = 144'hfb17fdb30203046dfeaffe19fc1201480182;
mem[516] = 144'hfc31fcf40086009200d5ff5dfd6cfdf3030b;
mem[517] = 144'h01be01e1fc4504d30166fcf70544fe08058c;
mem[518] = 144'hfdd5042807b6fd7efdda03bcfc5101d9fccd;
mem[519] = 144'hfe3e063b0d4dfa9a03260605014a0145f8ae;
mem[520] = 144'hfb24fdec0228ffd0fd5bfe55faff003e0134;
mem[521] = 144'hfd86ff9fff0501e4fe53fe33fa5ffc66ff84;
mem[522] = 144'hfb89fc47006903c5ffaafcb1fb05fe33fee0;
mem[523] = 144'hfc1301a809770281f9c40182fa9305c30287;
mem[524] = 144'h0066fd08fe9401d1010dfe3dfd03ff01ff5c;
mem[525] = 144'hfe90009ffe7dfe84fe4bff89ffc4009e00c2;
mem[526] = 144'hfbf2feeafb060263fef6feb4f9f0fdd5049a;
mem[527] = 144'hfbc5fbfeff7802dcfddbfd37fab9fcb700ee;
mem[528] = 144'hfc3dfb3cfcf200faffb2fc0b00c5ff53fcb0;
mem[529] = 144'hfd3cfb31000001fefed6fd1a0116019efe3a;
mem[530] = 144'hfbaef9a301bffbe0fa12faf00354fea401c6;
mem[531] = 144'hfe86fc1202aaff2ffc1afbf301c500e6fd2d;
mem[532] = 144'hffd5fc53fe54025d001cffcf024b01f0fd4c;
mem[533] = 144'h01c1fbbcf4450519057cff00007efbe8fe97;
mem[534] = 144'h00b1fff70020fbc7fe1304cf04d9035afe40;
mem[535] = 144'hff4301660154f8a0f96e054c03c302a00309;
mem[536] = 144'hfba4fd9b010d0055fe67fd3aff9e00ddfc7c;
mem[537] = 144'hfe38fd41fd9a0232fdf0fd3c034602a7fe60;
mem[538] = 144'hfdbcfb1ffdfcfe63fda6fbfe02b20086fd34;
mem[539] = 144'hfc58fd210120fa75fdd504740167fc63feaa;
mem[540] = 144'h002e01950113004d02a6ff06001600b10150;
mem[541] = 144'hfe5efe9bfec0fe2100f600030160fe9b01d0;
mem[542] = 144'hffbafe40002c06590073fc0502ce014ffdef;
mem[543] = 144'hff66fafd0091003dfcf3fae901cefe4cfec4;
mem[544] = 144'hfdacfe6cff3c00edffe0fe7bfdb5ff300138;
mem[545] = 144'hfeecfeb1feb1ff01ff78fe4ffec5fe2400ee;
mem[546] = 144'hffa4ffbfff63ff8a012c000bfe27fef9fe46;
mem[547] = 144'h0044006600dbff1bfe02ff21fde5fe96003c;
mem[548] = 144'hff4bff19ff2c00b3ffccfd9e00f7ff71ffb5;
mem[549] = 144'hff88ff83ff29ff0d00c00042fdbefed9ffb6;
mem[550] = 144'hfffcfe71ffb2ff53fda9fecefdc1ff290111;
mem[551] = 144'hfe70fe5dffd1009a002f00a5fdeeff3c00e4;
mem[552] = 144'h0069ff8dfffefef7ffeafecc008b0154005c;
mem[553] = 144'hfdddfe2c014bfde3ff32007b0136ffd4005a;
mem[554] = 144'hff3a00cc00ffffd3ff46ff670145ff9d000d;
mem[555] = 144'h00a3feefff6fff17003501b4fdfdfed8fffd;
mem[556] = 144'h004fff0bfe4aff07fe45fe4afedbfebb0008;
mem[557] = 144'hfeae006201640143fe4300d20070007a01bb;
mem[558] = 144'hfec00050ff3dfdf0fdacfef8ff62fdac00ac;
mem[559] = 144'hfe86fee1fe47fe8900580104febaff110122;
mem[560] = 144'h016dfcc9fb84ff33feb7fead05c200c1fe78;
mem[561] = 144'h000cfc9afddbffe4ff0dfe81056bff24fbd1;
mem[562] = 144'hfdc7fa89f70cfbf2026cfaa3023ffe85fed6;
mem[563] = 144'h0042ff3afde8fb46ffe2fec003defe75fe1d;
mem[564] = 144'h027ffc86fb59fb9e0039ff0a0210012ffc38;
mem[565] = 144'hffb8040afb08fc78029b00aa00d7fceff9e7;
mem[566] = 144'hfef5fd4bfa39fc770208007c040904480279;
mem[567] = 144'h0011f9b3f826003c01d0027d00b402a304ed;
mem[568] = 144'h007cff6afd6afd00ff77fe9e048fff5ffb7f;
mem[569] = 144'hff5900b8fe19feb202defe3a06f405a5fe6c;
mem[570] = 144'h00bafcccfe16fa8dffc9014f057d028b0070;
mem[571] = 144'hfe76ff87f9e202ab0362ffebfe79f975fab9;
mem[572] = 144'hfe47fd7a003f0065fff0004c0019019f0028;
mem[573] = 144'h00e8011cfec9ff1dff9aff5d00bffe77ff40;
mem[574] = 144'h0153ff3f000200f7ff19fe3501a8fefafc15;
mem[575] = 144'h003efc67fdbbfecaff90fd1a052900dafe0c;
mem[576] = 144'h01510191feb800aa0219ff1c0356040dfe27;
mem[577] = 144'h013fff48005bfe0201b7ff9504a802d2ff57;
mem[578] = 144'h036800dcfcf9fd390218031d0131fe0bfc1f;
mem[579] = 144'h002501abffe0ff14024bff5303a0ffa2fc90;
mem[580] = 144'h00e2fff6ffd6fefd0015001fffe702fcfd6e;
mem[581] = 144'hfe66ffc200d2f9ff0178002c010e00a90001;
mem[582] = 144'h019bffa6fbfc0142ff8dfdc10038ff42ffe4;
mem[583] = 144'h005d00b4fcf80140fff7ffeaff7bfe61fc75;
mem[584] = 144'hffebfeccff30015b0150febc02570239ff2a;
mem[585] = 144'h020a0241ff90fedc008b0033007a028dfdbf;
mem[586] = 144'h01970292fec6fee301a80009ff7b014700d1;
mem[587] = 144'hfd510383fc090126fd6ffc73010a0152fb75;
mem[588] = 144'hff3effce0099fff1fd3500f9fdf5fef60114;
mem[589] = 144'h013701a9ff070095ffc5feddfeb501730132;
mem[590] = 144'hfde200a301c4fed7039aff7102780268fd0a;
mem[591] = 144'h02c20062ffa0feb400b5fef200b701fafe08;
mem[592] = 144'hffdf00d00113fe420082ffeefde2fe85ffc3;
mem[593] = 144'hfe0f00e6015ffe4fffdb0116ff65016bfecc;
mem[594] = 144'h00d8ff9e0082ff0801f401b9fe58ff1e007a;
mem[595] = 144'h013e0167ffb1febfff2b00e5ff55ff4cfdce;
mem[596] = 144'hfdb8fe29006fff5cfe3ffe930145fe59fffc;
mem[597] = 144'h00c3ff7b017bfe36feccfef900c9ff920062;
mem[598] = 144'hff1fff6dff9c0092015a00f8fe53ff1800d0;
mem[599] = 144'hff5e0096fe9cfe41ffffff2efe46feb6014a;
mem[600] = 144'hfedafe7afe73ff1200030073fff7ffa0fe5d;
mem[601] = 144'h012f0088fffb004d00210010ff64ffe1fef6;
mem[602] = 144'hfea8013e00260041ff56fdcf016dff96ff21;
mem[603] = 144'h01cb0019ff55feaaffc4ff2700e601b70177;
mem[604] = 144'h0177ffad0064ffd400700080010201d401c4;
mem[605] = 144'hff99019d01e0013b01a900b0012e00ec0007;
mem[606] = 144'h00e7fed0ff04fe4ffdf00149003efefffdba;
mem[607] = 144'hfea2fed4fdd0ffff00f20129fe3f001a0175;
mem[608] = 144'hfbcfff780056008a0084fe9400acfe0afde0;
mem[609] = 144'hfeb4008f016afe6cfdf0007afff9fec9fda8;
mem[610] = 144'h005cfd5affddfe56fe79fcb9007bfef903cc;
mem[611] = 144'hfbd5fe230161fffa014aff8cffb7ff93fe92;
mem[612] = 144'h0071fe9f01a0fea300c9012f01710021fe20;
mem[613] = 144'h00bdf9d3ff1c05b7ffd2ff7efc2ffad4fbd6;
mem[614] = 144'h00df00d701f7ff2dffe4012e03cd023b0063;
mem[615] = 144'h00f1ffc403baff58ffb40127025a03ae0314;
mem[616] = 144'hfc16fdcefe82fd6c0142fe9dff8afec9008c;
mem[617] = 144'h00ecfd99fefc001bfe1801f4052d004cfef3;
mem[618] = 144'hfe55ffd9016a0092007a00c1011f02830063;
mem[619] = 144'hfe73fc26026fffd301b00312fdf8f977fd90;
mem[620] = 144'h00aaffcf01ddfe92fecfffb10039009f0036;
mem[621] = 144'hff17005700d300cc0126ffcaffa801820002;
mem[622] = 144'hfc83ff4600ebff1dfc9ffdd802b402d100e0;
mem[623] = 144'hffc5fe130000fd8aff5aff380261ff5a00ff;
mem[624] = 144'hfecbfddcffd6ff73008bfe5bff81ff6dfef2;
mem[625] = 144'h0019013dff31016901a9ff4601210110fe7e;
mem[626] = 144'hff9fffb6fef9fed3ffc500aa006f01c001b7;
mem[627] = 144'h0107000efedffff500650033ff16fef300e8;
mem[628] = 144'h0186ff43ff90fe880185fedaff78001a0052;
mem[629] = 144'h0064ff9aff20ff8bfee3005c010f009ffe47;
mem[630] = 144'hfe2e00fe0184002dfe3300d60044018ffe8b;
mem[631] = 144'h0096016dfe3cfff0ff69006501bb00f3fff8;
mem[632] = 144'h00acff3fffaafeadfebb0131005dffa9fe0c;
mem[633] = 144'h016d00c4feb0fe6afe03fdd2008eff86fe02;
mem[634] = 144'hfdddffdcff91ff79ff04fffa0132014cfe86;
mem[635] = 144'hff270194ffad01960037fd8b00d80115ff98;
mem[636] = 144'hff3201cdff4dfee8fed8fe8dff7101c301bd;
mem[637] = 144'hff47feafffa2006c00f3011e01d9fe41009e;
mem[638] = 144'hff7300d7ffc0019f0023ff9001750161ff67;
mem[639] = 144'hfeb5fe38ff6efeb8ff550161fe2b0013011c;
mem[640] = 144'h01fffc3f0006fd47ff7c006207ad0271ffc7;
mem[641] = 144'h00e0fddafd310017fe7c00cc0a4001e00099;
mem[642] = 144'h0269ff6800d2fe11008a08e904b602c7037d;
mem[643] = 144'h003a011b0157fe1600fb059105f103040176;
mem[644] = 144'h04a80023fed2ff50010c026a058c038e01ed;
mem[645] = 144'hfe5cfb50f5f103f1ff3901befdbaffecfe02;
mem[646] = 144'h0565016f00a0007503ea06d005de050a022f;
mem[647] = 144'h019c02290181ff1c08ca078500f2041f0471;
mem[648] = 144'h00a2fdddfe73ffa2014d0326068e01d30162;
mem[649] = 144'h04ecfe2cfeac0396009301fc08bf04b6ff64;
mem[650] = 144'h03fe019dff40ffddfe63019d071706680026;
mem[651] = 144'hfc68fe99fe53fa0ffd2ffaa0024ef9f7012e;
mem[652] = 144'hfea1fd230088fef9fdf4fe88ff3902460033;
mem[653] = 144'hffc50011fee5ffc90090ff4700d50038013a;
mem[654] = 144'hfb48010a01810116fdf5003d06b1fd83fcb4;
mem[655] = 144'hffc7fd87ffd9ff9100af0043075d0160ffa4;
mem[656] = 144'h0155ff700003fe330009febb001afe8a0093;
mem[657] = 144'h00c10044014bfee9001dfe3b0073fddeff35;
mem[658] = 144'h005c00bffe74fe1100030122ff980158004a;
mem[659] = 144'hff7f015cfdfe012bff1dff2e0108ffe30063;
mem[660] = 144'h00a8ffc3006effe9ffea007bfde7fda7ff9b;
mem[661] = 144'hff78fef8fdebfdcf00690030ffc50115fe79;
mem[662] = 144'h003d0133fee10185014cfe09fe38fecbfe47;
mem[663] = 144'hfdc1fe0900860084fdeaff1f009f011dfee6;
mem[664] = 144'hff68000100a300e100dc00580048ff47fe13;
mem[665] = 144'h0076fdbdff0100defebcfdc6fe3001c10049;
mem[666] = 144'h00ba0139fdfe00a3fe9e0017fff1fe6cfeaf;
mem[667] = 144'hff32fe8d015e009eff240023014f01160088;
mem[668] = 144'hff6bfedb016f0109fe9a007101b9003ffe5e;
mem[669] = 144'hff7a00a200aefe3e000601ca01ccfebfff04;
mem[670] = 144'hfeb400090098ffc9ff1cffa10160014a0061;
mem[671] = 144'hfe05fe23fe7800e5ffb0fefb0063ff9afe0e;
mem[672] = 144'h0255fda3fd4afd2e030d030e0019fc59fad5;
mem[673] = 144'h0343fce1fdcafcc005a40120009afb95fab2;
mem[674] = 144'hfd9ffc5ffb8206730516fbaefc60fd65034c;
mem[675] = 144'h0128fe2cfbe60212034400c8011afb4fff36;
mem[676] = 144'h0239fe09fc0f012103cb02490381fd4cfe92;
mem[677] = 144'h005003e90321f9ab010b02a9ffb2fc16f748;
mem[678] = 144'h020bfcb4fe2f037603fc0241007500fb02a4;
mem[679] = 144'h002bfd6000b00b5efe7bfeaeff4b05be0828;
mem[680] = 144'h02830001fc7600560389ffa2ff59fcaefe7a;
mem[681] = 144'h0122ff9afcccfc910522fffe0572ffd0fb84;
mem[682] = 144'h021efac5fd21fdf3055b03910216fd9bfc35;
mem[683] = 144'hfd74fdcff96d09db00bf0050fa92fa2afd9d;
mem[684] = 144'hfd51fd70002000f8fe83fdffff5600630091;
mem[685] = 144'hfe8aff2400f2006f0144ffcbfe59fec4ffa4;
mem[686] = 144'h038205ccfed1fbad024f00c101b0fc0bfbdc;
mem[687] = 144'h00e9fccdfa7100ae044200970363fb7afc69;
mem[688] = 144'h013601da0425023aff47fc36ff30ffbc0361;
mem[689] = 144'hfe9b0013016805050152ff7d000eff1c02d2;
mem[690] = 144'hfe54009f03a40028fecf04c902ceff4bfed5;
mem[691] = 144'hfe8cff5104910547fe2afe0b015d02ff030e;
mem[692] = 144'h01f50017033e03b8fd49003c0221ff0dffe8;
mem[693] = 144'h00aeffb8f7ed0564010f0035049d029bfb17;
mem[694] = 144'hff7402a705cbfd9cfcd0ff7102a9fefefcbd;
mem[695] = 144'h008bffcd05e7fbbf0033039c017d0093fc9a;
mem[696] = 144'hff620073050a0429fe52fdea01cc021d0154;
mem[697] = 144'h016804f101b10160fc8ffe70ff7bfea30025;
mem[698] = 144'h023c027902890574ff55fe9f0046001d00ab;
mem[699] = 144'h00f4ffb80301f951fb080178006c028d03e6;
mem[700] = 144'h00b3fe5dfe88fdaa01f80179005dff7a00e4;
mem[701] = 144'hffb90021fe6d0160fe7c012e0100ffc2010c;
mem[702] = 144'hfd7efd7d0121071100a1ffabfd8d020c03f3;
mem[703] = 144'hff4dff0203e20566ff67fdd1021e007202ad;
mem[704] = 144'h028700f105bd04b40170feac02cefd5d01fa;
mem[705] = 144'h02b2023b0552042f01e9fef3ff50003d00fa;
mem[706] = 144'h046bfe07fb6cff72fcbbff4100d4faa4ff97;
mem[707] = 144'h01d9036b02230402fef3fc8902a90119008a;
mem[708] = 144'h00bc031401b8022700e4fd250180fd7e008b;
mem[709] = 144'hfd72fb13f64dfa650237fed5fd37fa8cf4f9;
mem[710] = 144'h0183008600cfff8efebafce2fe49fbcc0155;
mem[711] = 144'h00d9faebfd65f9b3faad01fffffefc53fe13;
mem[712] = 144'h014f01cc051104e4027ffcc3013100a40152;
mem[713] = 144'h00a6016a0331031d00edfcdbffd1fed4fcfa;
mem[714] = 144'h01d60241053c054103580005014900affe0c;
mem[715] = 144'h023ffdf5f783f7b6f876fe5d010dff95fb7c;
mem[716] = 144'hffbafec3ff6dfe1dffae00ebff11015302ae;
mem[717] = 144'h0019fed3fefbfe930020ff38ffef018dfe8f;
mem[718] = 144'hfdf9023505690412048dffc1019002ee0234;
mem[719] = 144'h02990163045005b002b8ff9a01590002ff65;
mem[720] = 144'hfc38fd04ffe3009bfd48fd1f016a0154ff55;
mem[721] = 144'hfe34fb640013ffd1fd5cfd4500a3003fff73;
mem[722] = 144'hffb2001f06c0fc58fb7f00c302ab0437ffa4;
mem[723] = 144'hfdd1fdb702c1fddffc2400a1017d04c50174;
mem[724] = 144'h00ddff9fffc2006bfe65018f01f00142ff5b;
mem[725] = 144'h0234fd23fe4906f7fe8bfe7a00e103a608f7;
mem[726] = 144'h02db034e025bfbacff860390035c0200fb6e;
mem[727] = 144'h00ce075a049ffa49ffa403cf032403f00085;
mem[728] = 144'hfefffebcfea4ff5afcfbffab016d03820029;
mem[729] = 144'h020cff87fe81028bfba9fed6ffb8ff59fef4;
mem[730] = 144'hfd1cfeaa009e010bfe29000f014001acfed6;
mem[731] = 144'hfdf2fc36076ffe000186fffd0248fddb04e7;
mem[732] = 144'hffdd02b100ddff4c02edffc4feed00d9025a;
mem[733] = 144'hfe60ff0d0000ffe3feacfead015b00e1ffbf;
mem[734] = 144'hfecafc71fc530153fd37fc5000c8ff660101;
mem[735] = 144'hffaefef2ff4f014cfbf6fd7000b301f80161;
mem[736] = 144'hfe1f0063fea2fec1fe3f00d4fe94fef50053;
mem[737] = 144'hfe3e0149fe96fe25ffd9fe70017cfdf1011b;
mem[738] = 144'hfe68ff2c000efeba0146fecdfe58fe3cff35;
mem[739] = 144'h0015fdd0fdbe003a00a100bd010efe33012b;
mem[740] = 144'h007afdd2fde10105ffecff5b00dd00470101;
mem[741] = 144'hffb20022fee3fdcffdcc0140fe4ffe730096;
mem[742] = 144'h00c1fdc2ff72003efdeb017f0090ff67fece;
mem[743] = 144'hffbbff43002101bdfe82ffbe0001ff1c012c;
mem[744] = 144'h00960051fe57ff70fdd4ffa1fed800f8006e;
mem[745] = 144'hff54fea001d2ffc90048fe2c01b701440025;
mem[746] = 144'h0009fe33feca015d0056fe2efeb101490107;
mem[747] = 144'h005700f100d4009b00910043fe7b00f30179;
mem[748] = 144'hff8700ff012501be00a9fe23ff57fe4fffe7;
mem[749] = 144'h0055fe8afff801c0ff940078011afe2600ed;
mem[750] = 144'hfe99fe17fe45fef8feaffef0ff94ffc1017c;
mem[751] = 144'hfef8ff91ff2000b5fe99006fff84016efdce;
mem[752] = 144'hfe51fe2c028000a5ffc8fef507200512ff41;
mem[753] = 144'hff7dfcd8009f03a80023007506ec0496ff9b;
mem[754] = 144'h0036036707bafb5afe7405da066c0397ffa6;
mem[755] = 144'hfd99fff703d000c60071049103f405cf00b2;
mem[756] = 144'h024fff53037202c4fef2022304be03f70015;
mem[757] = 144'hfd93f85df69604d1fc2c0228ffa2016a00bd;
mem[758] = 144'h033604500696035105d808b105df0341fd42;
mem[759] = 144'h031509b103affb38042c037602be0235fca9;
mem[760] = 144'hfcb1ff190157023c0020ffbc063904c50027;
mem[761] = 144'h02a0fd5f00b502a8ff9402db075605c9fe6e;
mem[762] = 144'h0404012303bf04f1018402d7078b04e501d9;
mem[763] = 144'hfb99fccf0101f3d1f8eefbf10461fd2e0341;
mem[764] = 144'h0002fef300db00b60117feeeff6e0049ffe1;
mem[765] = 144'h020000ce00df01b7feda00fb011300c9015d;
mem[766] = 144'hfa7bfbd60088004e006cfe93048801680231;
mem[767] = 144'hfddcfdf50292010cfeff027803c501b3ffea;
mem[768] = 144'h010103de0092fc7c024c03e3ff1400e7032a;
mem[769] = 144'h00b400200083fe3300f703cafdbc00e902e7;
mem[770] = 144'h02d4078206a809c204f90c9e01740236fff5;
mem[771] = 144'hffd903bf009a051a023b0555ff69ff9d0240;
mem[772] = 144'h00e10285ff5401fd0284048cff1500d30228;
mem[773] = 144'h00cd0293091e0324fe62fe4201160740050f;
mem[774] = 144'h022102f1054e04dd010f04a20019fe36fdfb;
mem[775] = 144'h0241046b06e6065006e501da00f4014dfdf3;
mem[776] = 144'h017900c60096021601be0353ff36016a0377;
mem[777] = 144'h029401f6ff7dfda2fdec0319fde3fcfcfe95;
mem[778] = 144'h034301f2018c02ea002b01acfcc600c7ff6c;
mem[779] = 144'h01d1006504b008cbfe9efcd6005b0313082d;
mem[780] = 144'h008bff0eff260038fe70fff900c2011000a4;
mem[781] = 144'hff4fff0700fcfe91ff1601deff11fe7fff91;
mem[782] = 144'hfdae00aefa9afc71010c061fff68fce80041;
mem[783] = 144'h005501150009001602c4061c01a301130196;
mem[784] = 144'h0098ffad0386044601d1fcc504f5027002ba;
mem[785] = 144'h000b009604e403b5ffcafcd701b3ffe10281;
mem[786] = 144'hfec2ff4200affac4fa3f0179042e003701da;
mem[787] = 144'h00dc010705ef0281fca600120206035600e2;
mem[788] = 144'h0233ff250490016bfd93ff7d00c60042008d;
mem[789] = 144'h0100fa4af5e605a102deffb4ff18fe53f8d3;
mem[790] = 144'h02b4016f04b6012aff45ff1e0527003a013d;
mem[791] = 144'h025d01aa0021f855017d070c046b018c0073;
mem[792] = 144'hfe3900f40497042a0002fbb9033a02f50274;
mem[793] = 144'h02ea0180035a0432ffd4fe99032afee4020d;
mem[794] = 144'h030b00a004a703f20016fdb604ff0190ffc1;
mem[795] = 144'h00edfd3f011cf3caf78504b8ffa40067ff84;
mem[796] = 144'hfde600f3ff4afe2cffa8ff08ff82024d0218;
mem[797] = 144'hfeb3fefefede019cfe710044ffe8ffe6008b;
mem[798] = 144'hfd06fde203b405a7fdcdfbaf03a9012701e7;
mem[799] = 144'h0168fd9405fa0446fe5efd6703af0320025b;
mem[800] = 144'hfd86feb0009a01050199fefffd68fe450091;
mem[801] = 144'hfe9900c9feeaffdc00ebfdccfebe00c1ffe6;
mem[802] = 144'h0002013ffdc0fff2fdf6fefafe72ffb2ff55;
mem[803] = 144'hff8e00aaff5000a3ff57fddeff6e0072ff41;
mem[804] = 144'h00bfff9e00b10007fe220139ff3e005d00e0;
mem[805] = 144'hfd9efeb3fe83fec4017eff1cfeecfee9fdb6;
mem[806] = 144'hffffffbdff21fe15ffa8ff9aff65fda6ff41;
mem[807] = 144'h00ea0036fdb3ff54feceff4fff06fe0bfde8;
mem[808] = 144'hfe06003d0053fe9b008afe7a00faffd4ff3e;
mem[809] = 144'h0091fe900064fdfb0197ff38fe170140fea3;
mem[810] = 144'hfeb1ff61ffb700b9ff9a00ebff2ffd35fef1;
mem[811] = 144'hfed60145fed1fdd4ffd8fdd0fd86fe96feda;
mem[812] = 144'h00c5008b018affca018cff77006401c7ffa1;
mem[813] = 144'hff38feacfeac01dd005e01900102fe86ff4e;
mem[814] = 144'hfda1ff17ff95fffafdadfe73fff500610134;
mem[815] = 144'h002dfd71008ffe83febffe28fee4fdd9ffc4;
mem[816] = 144'hfdd4fccbfd23ffae030d0218023afe49fce2;
mem[817] = 144'hffc7facafac1006a03e901b9ffc6fe76ff45;
mem[818] = 144'hfdf2fb260268057f0088f9e20275fd010450;
mem[819] = 144'hff17fbc0fc890116015402e80078ff4d016b;
mem[820] = 144'h02cafebefd59fefb010900bf041500b1fff8;
mem[821] = 144'h02de07abfb78fea40172041b003cffcff770;
mem[822] = 144'hfe64ff6b0106009d038bfe21044d03ff063b;
mem[823] = 144'h029cff8c044301befdddfb7d046701e40723;
mem[824] = 144'h0048fddafbdc0076040f02abfee5fe8dff44;
mem[825] = 144'hff48fd2ffbfe00fb04ad02360446016d0050;
mem[826] = 144'hfebefac0fc1dfd7700a802be01bcffadfe97;
mem[827] = 144'hffddfd430262042c02440151fd9ffc110192;
mem[828] = 144'h008affc80156ff3effed015cfd03fe2dffbe;
mem[829] = 144'hfe8fff71ff96007f0101ff840180ff94ff0b;
mem[830] = 144'h027cfe26fe4f001201f4031202dffe7bfb6e;
mem[831] = 144'hfdacfdfefbc2fe50013d03cdfff6ff2ffd6d;
mem[832] = 144'hfd1e04d401fafff1fe90ff70f859009201c7;
mem[833] = 144'hff1d03420084ffa7fec001a6fac200e600c3;
mem[834] = 144'hfbb3041d0135fec6ff6ef97dfe44ff2bfda9;
mem[835] = 144'hfedaff7dff3dfeb3fef2fdcdfa32fe66ff50;
mem[836] = 144'hfc3f0324033d01aaff88fe26fcdffe5b0075;
mem[837] = 144'h00880a8e0ce0ffb8ff5702b8048105b00af3;
mem[838] = 144'hfb1802c3019ffde1fbfffaa0fdddfb54fd34;
mem[839] = 144'hfb08ffe7011bfef3f97af9de01dbf921f83d;
mem[840] = 144'hfdeb03a70010ff4dfe630008fb0101ad015d;
mem[841] = 144'hfb08042efe73fec9fc53015bf8b1fd11035d;
mem[842] = 144'hfa4202fa01a20106fd21fd01fae3fee9ffaf;
mem[843] = 144'h021e07ea0589037106a10283ff28086803e3;
mem[844] = 144'hfff6ffe0fecc00c800f3016fffe1ff7cff97;
mem[845] = 144'hff8cfea6fefafe2800290178fe9affb701d0;
mem[846] = 144'h023e02280074021e018a028bfb99019c035c;
mem[847] = 144'h00200415026d01f4004efe40fc59009202b7;
mem[848] = 144'hffb4fc4cfe23fc62ff6d042efd0a01f60424;
mem[849] = 144'hfd8dfc3dfb2afb97feaa04e7012001430320;
mem[850] = 144'hffee01f901d7054b0563fdfefdde025c0456;
mem[851] = 144'h0064feaef96f001202ce0259ff7302cb031d;
mem[852] = 144'h002dfc5efd6cff30000803c2fe64027d036f;
mem[853] = 144'h011707630e5c0125ff9a033f0157ff8801d2;
mem[854] = 144'h008fff0ffe0d039201ff0242fed805460452;
mem[855] = 144'h02dd039707d80a20051dfd930190029f038f;
mem[856] = 144'hff2cfd9ffb6ffe60006d0378016502b90382;
mem[857] = 144'h0088fd5cfbf4fafd00b50330005b02480514;
mem[858] = 144'hfd51fdaafcf5fc32033d0684fee5004a02fc;
mem[859] = 144'h011602fe01c8083208b90491001301e8ff33;
mem[860] = 144'h020a007a018d0205fd19fe6ffef1fdf7fcb0;
mem[861] = 144'h0174ffeffe96ff96ff710077ffde0197017c;
mem[862] = 144'h018c0017fc80f6f3fd7a023eff51fe2bfeba;
mem[863] = 144'hfe65fea5fd7cfb3c01da043dfe64000b0308;
mem[864] = 144'h03ce0431fdcdfb0afe180391017801330489;
mem[865] = 144'h01f10434feacfa05ff8601f90270024f0359;
mem[866] = 144'h053a04c5fcec04ca0366096801bb01e00340;
mem[867] = 144'h00f60488fbaefd9a007105b60196021a034d;
mem[868] = 144'h02dc00a8fcffff4f01b1034b01f90358022d;
mem[869] = 144'hff92042b0c280335fc89fcec000e03a501bf;
mem[870] = 144'h04eb0185f8a201bc03600170fe6f019104ea;
mem[871] = 144'h03980013fb330415071b00a5fdf8010f02cb;
mem[872] = 144'h04b10341fcaefaed0164042a025802710137;
mem[873] = 144'h0295ff670011fca3fd7e034901acfff001f7;
mem[874] = 144'h037700520123fd1efe66010c03670045060b;
mem[875] = 144'h0209025afeab0a8304d4031a02470175013e;
mem[876] = 144'hff5d01c20177ff22fd2dff6701a8004e0055;
mem[877] = 144'h01a20145ff590036fe8000f101b3001c0165;
mem[878] = 144'hfd17011e01b5f7a8faea0143035e006d0126;
mem[879] = 144'h01140331fe7afdfcfff503ef0180034b041f;
mem[880] = 144'h03c1fe32fed0fd2b010dfed805e201300156;
mem[881] = 144'h038601ab009bfcfdff64fe53047701ff01a8;
mem[882] = 144'h01f7ff2bffbf02520345040101990252039e;
mem[883] = 144'h0206009eff54ffbb02ea0008030d020001c3;
mem[884] = 144'h02f0fecb00d1ffbf022afeb303cf024c0319;
mem[885] = 144'h0046fa5dfe790163fd70fd3ffc2afeb2fa99;
mem[886] = 144'h03bdfea3ff4a01cb01aa003103590416031c;
mem[887] = 144'hffba000dff7c04f404930243fead0171059c;
mem[888] = 144'h03490132017eff40ff6001dc0316019d01b8;
mem[889] = 144'h032dfdecff590055ff5efeb3040c012d003c;
mem[890] = 144'h05ddfee7ff58ff6e023a017804460398048e;
mem[891] = 144'hfd15fc1cfd8e028bfbaafc92fee2fe3cfe7a;
mem[892] = 144'hff46ff330004feb5ffce0026ff3c028a006e;
mem[893] = 144'h00e30013006601dd006e01250137006dfe93;
mem[894] = 144'hfdbffdab0018fd80fdef00e70237fe74fe30;
mem[895] = 144'h0155ff380020fec400dafecc060502f80372;
mem[896] = 144'hfc5ffcecfbdbffaafd80f88efb87002b003d;
mem[897] = 144'hff3dfc42fcdaffe6fcdef91cfbe70046ffe5;
mem[898] = 144'hfd67fe1e06ac0211fd46f84efc83ff9800d0;
mem[899] = 144'hfd39fc55fedcfefffd6df7f5fcea005500ae;
mem[900] = 144'hffad00b000e9fe81fdb6fc0cfe570077ff26;
mem[901] = 144'h02290752021f07cb02f0fea400b700330557;
mem[902] = 144'hfdb302b40566fff9fb29fcc1009802a7ffde;
mem[903] = 144'h025a03f10c5400a9fb8602b001fe047f01e9;
mem[904] = 144'hfcaefc5afc06fd33fd5cf8befc24fff901fe;
mem[905] = 144'hffadfe87fcfaff9cfbe5f9e6fe67ffa2007d;
mem[906] = 144'hfea7ff0e0027fddefeacf7b7ff8500abfff6;
mem[907] = 144'h001d01f705f303a104020534023603cdfe12;
mem[908] = 144'h015200a7fff800ac02db0085fce80132ff93;
mem[909] = 144'h002ffeaf0077fec4ffd80107019dfec9018c;
mem[910] = 144'hff77fffafa130118fea1fad8fef303ed034c;
mem[911] = 144'hff87fe13fe92fda0fdf0faedfd1d01d3ff4f;
mem[912] = 144'h004efd85ff63feeefd75fdc4ff02ff4dff0b;
mem[913] = 144'hff7bfffbfe0600e5fff500e8fe8ffe5bffea;
mem[914] = 144'h00effe8cfee7002afffffd7afe43ff57fdb4;
mem[915] = 144'h0016ff12fe7f003ffd74fe3aff400057fe81;
mem[916] = 144'hfe37012fffaeff0a010bfe3f007900fbfe0e;
mem[917] = 144'hfe43fe430080ff8cfe71fe20fe81ffc1feac;
mem[918] = 144'h00120102ffbbfeb200570019ffc8fdd5fe72;
mem[919] = 144'hfe87ffcf0053fd89fe87012b000d0006ff64;
mem[920] = 144'h00cdfdcbff5dfd6ffe19fed1fd80ff23fde4;
mem[921] = 144'hffeafdb0ff1dff19fd9500acfe46ffd8fd75;
mem[922] = 144'hff5cfe75ffb0fe3dff97ffa70095feab00a2;
mem[923] = 144'hfffaff82fed90033fe33ff1afdbeff0afe82;
mem[924] = 144'h012200f9ffc3ff8100bb0061fee30008005d;
mem[925] = 144'h0076ff50ff3a01bf010d018d0121018601de;
mem[926] = 144'h006500bcff53fe9cfe90fe1a004200d4fe7f;
mem[927] = 144'h009800e30038ff8d00d8feb1ff29fee5fea7;
mem[928] = 144'h00e304ed0095016e025effbbf9f500d50106;
mem[929] = 144'h010804ed00bf027801300086fbaa01810250;
mem[930] = 144'h02610612023c017bfb63fd7200640012fac0;
mem[931] = 144'h0066029c02bb02f4fe50fc63fd1002b8fd99;
mem[932] = 144'hfd0a04740261024cff02fefefcdcfe0cfdc9;
mem[933] = 144'hfeacfc0103b6fc410208ff39023a053d0609;
mem[934] = 144'hff4402ad0350017afd33fdd5fed4fc02fb14;
mem[935] = 144'hff330176ff16fcb9f933fdaf00e6fb7ff51d;
mem[936] = 144'h004f012000e1035b000afea0fcb202aaffba;
mem[937] = 144'hfc5001e102b0ff13009efcf7fa62fc5effe1;
mem[938] = 144'hfcbe02fb014f01320035fe3bf988fe7cfe6c;
mem[939] = 144'h019b021fff37feacfb6bfd5001420415ff6a;
mem[940] = 144'hffe3ff56ff4a004d00ceff56fe28fd43fec0;
mem[941] = 144'hfe1aff3cffe900de01450140fe8f0153ff31;
mem[942] = 144'h0176fdf300a60182037b025bfadd01e702e2;
mem[943] = 144'hfe1204c8014900fe009cfee1fb9f024f005d;
mem[944] = 144'hfebafe3cfef0fe31008cfe5b011c0151ffcf;
mem[945] = 144'hfe88012d0076feb2ffcefdcffdfaff19fe92;
mem[946] = 144'h0046fdb2fd88004efeacfef00025008afe11;
mem[947] = 144'hfe7dffe500c1fe59fdcc00c2fdadff66ff40;
mem[948] = 144'hfe46ffafff4b0050fd910114fdb8005800d9;
mem[949] = 144'hfdfbfea4ff01fd9efe6bfefcfe7a012bfded;
mem[950] = 144'hffabfe07fde20007fdef005ffeb20131ff6f;
mem[951] = 144'hfdd100dffde6ff2f00f8ffe9ffafff8bfdcd;
mem[952] = 144'hfd74ff62fe2fff8cfe30fda2fe17009c00c6;
mem[953] = 144'hfd9efe4b00f400e5fde7ff64013000ee0068;
mem[954] = 144'hfff4fe89fed6ff39fe3f007b009ffe4cff52;
mem[955] = 144'hff79ff82fe77fd5f0109ff0e011ffe45009e;
mem[956] = 144'h008b011a00d1002200b4ff5fff0cfe88016a;
mem[957] = 144'hff2201cdfeeb004affd20177018e01d6019a;
mem[958] = 144'hfe4efe50010fff94fd7b00ddfd93006dff39;
mem[959] = 144'h003700beff2cff3fff03feadfe67ff4cfeb0;
mem[960] = 144'hfefbfe2b00780105ff53fe38fe09ffe9fe75;
mem[961] = 144'hfe8aff1500f0ff1dff9cfef50168ff27ffa0;
mem[962] = 144'h01c70049013c0178fe2400ce0141ffd2ffbb;
mem[963] = 144'hff9cffa7fe8400bafef9fdc6ff8bffaafdff;
mem[964] = 144'hffdf001fff7afdeefeadff58005fff0f00b0;
mem[965] = 144'hff0bff16fef5feb1017e0129fdf9ff27016f;
mem[966] = 144'h002f003a006afddbfe8400e3ffe6fe61ff9e;
mem[967] = 144'hfe990098fe7effe50045ff70ff4dff34004c;
mem[968] = 144'hfe3100f2fe83010d0054ff54fe0aff7afdfc;
mem[969] = 144'h0096ff960013ff0aff4d0086ff8e0138ff50;
mem[970] = 144'hffb9ff160085ffebffd000ee007eff5e014c;
mem[971] = 144'hff57fe4aff35fdd8fed7feb90117feb4ff47;
mem[972] = 144'h0044ffecfe40ffdc014aff65019100b800cf;
mem[973] = 144'hff19ffd8fe8900b0005201c300480109011e;
mem[974] = 144'h0123fe61fe91febf0094001afdff001efe37;
mem[975] = 144'hfe5cff3cffafffc10029ffcbfdfafee4fe7a;
mem[976] = 144'hfff600c3ff78fdf6fd40ffbefe62ff59ff31;
mem[977] = 144'hff34ff94fd8afec2ffbdfcd9ff88fd3dff59;
mem[978] = 144'h028f00defdbc027affd8fd860033fd51ffef;
mem[979] = 144'hfe2f00aefddfff0dff84ff97ff60fceffd8b;
mem[980] = 144'h0076000e0201fd8afe46ff7dfeb3ff5bff29;
mem[981] = 144'hfefefdec0349fffffe37ff99fedffdadfe05;
mem[982] = 144'hfea702a30247021bfe730031004f0007fe62;
mem[983] = 144'hfe1bffa2ff10033cfe56fddafe25ffb8ff45;
mem[984] = 144'hff9b016efe460000fe12ff66ff30fe6a002b;
mem[985] = 144'h011fffd9005cfd6afe9701dafe24ff20fda2;
mem[986] = 144'hfede00a100b7feefffaafd08fe04ffb2fe1b;
mem[987] = 144'hfcfdffe5fea7ff9cffb50058fe26fe5efe7f;
mem[988] = 144'hfff901c2fe6b0011ffa401d700f4014500ac;
mem[989] = 144'h01cdff1f004afe61ff000198ff8100c9feec;
mem[990] = 144'h01f7fce9fd14fd2a02baff8effeaffd4001a;
mem[991] = 144'hfff50253ff7efe50ff24fea2fd5cfcd4ff85;
mem[992] = 144'h03fd013e02a5036fffc8ff7803befde3fedf;
mem[993] = 144'h016502cc03ae04f6010101dd03cc009d0151;
mem[994] = 144'h01e6fe240279fe8bfd5e06c3ffc4ffd004fa;
mem[995] = 144'h033502d701850372fefc00b50051011802fd;
mem[996] = 144'h018b027801fe0303002101b4031d01350175;
mem[997] = 144'h014dfd18f4a7019d0014fe2c00530007f6c7;
mem[998] = 144'h01e400640098003801a800be01f7010200b0;
mem[999] = 144'h0364febaff44feec054d059eff9202ed0308;
mem[1000] = 144'h03ed023e023902b5ff5e00d000dafef5ffb2;
mem[1001] = 144'h04400170017b02d0025800c801ddfccfff55;
mem[1002] = 144'h05a801530242068d00af002d02cb00bb0156;
mem[1003] = 144'h0236ff4b0273f60af6beff3bfe66fd8b0672;
mem[1004] = 144'h0055ff41009a00c6020cff6401b3025cff7b;
mem[1005] = 144'hfee8009b0003ffc800d00116fff1fef6ffc1;
mem[1006] = 144'h012601d004fc04c701f2014603adfd14fed1;
mem[1007] = 144'h010e013a04ee045501e3015c040e006500f2;
mem[1008] = 144'hfed60097fd47ff660257018bfff1fe93fe03;
mem[1009] = 144'h00d9ff39ff1d005702c5fe48008ffd25fc66;
mem[1010] = 144'hfd22fbe4fcb205ea01e60024ff90feb800f4;
mem[1011] = 144'h0051fdfdfdc1ff190157fd64fea7ff8f0047;
mem[1012] = 144'h00b4ffaafd9d001a01d2fe7cfe8cffd30000;
mem[1013] = 144'h0228fec7fd2701cc03b50323ff9ffcf8f83a;
mem[1014] = 144'hff5efd37ff840284fe6601c300150047018f;
mem[1015] = 144'hfdf7fd67057a0845fc0201c80137048c0785;
mem[1016] = 144'hfe66ff15fd59fed400b9fde3fd88fbe5fd08;
mem[1017] = 144'hff1dfe36000ffd2e01f9feb5019afd14fca5;
mem[1018] = 144'hfe0d0065feca002e014600f700fafea60000;
mem[1019] = 144'hff9efe70fa7609f5055d01f4feabfb4dfc2e;
mem[1020] = 144'hff2d001a01a8ffa1ff40017fff0efe97ffb8;
mem[1021] = 144'h005afe30009dfe3cfee3fe25fead01ba007a;
mem[1022] = 144'h013a004d0028fea90095ffbaffd30035fcd2;
mem[1023] = 144'hff000022ff4efe5a02c6ff0efe12fc25fe4e;
end

always @ (posedge clk) begin
	q_a <= mem[addr_a];
end

always @ (posedge clk) begin
	q_b <= mem[addr_b];
end

endmodule