`timescale 1ns/1ns

module wt_mem1 #(parameter ADDR_WIDTH = 11, DATA_WIDTH = 144, DEPTH = 76) (
input wire clk,
input wire [ADDR_WIDTH-1:0] addr_a, 
input wire [ADDR_WIDTH-1:0] addr_b, 
output reg [DATA_WIDTH-1:0] q_a,
output reg [DATA_WIDTH-1:0] q_b
);

reg [DATA_WIDTH-1:0] mem [0:DEPTH-1];

initial begin
mem[0] = 144'hfbad005b1176ebad01041380f8cb136c1fd3;
mem[1] = 144'h167e00220f3210011cb7f50a14581dd01959;
mem[2] = 144'h02da04affb46007bfff8f8c400510143f7c8;
mem[3] = 144'h07f006b500b304a60a8c009dfee2ff4a07bf;
mem[4] = 144'h05cb03c6019a0bdb095af8b1ff9bfc9cf65b;
mem[5] = 144'hfe6608b0077f0655052903b4fe79034700b8;
mem[6] = 144'h09e8fd5df30a05edfe00f01dff02f098f653;
mem[7] = 144'h024706b1032a07c7022c0911006c02be0315;
mem[8] = 144'hf3c6ff500c3302da05a209a904fe0285fe4a;
mem[9] = 144'hfb99f64d035701cb0798ffce09e403bc03d1;
mem[10] = 144'hf2940b0a0f6bfe6f0e5a0ea70f620eaa0b7a;
mem[11] = 144'hf2a3f97503f7f5b0fd3e096cfee2069f0b52;
mem[12] = 144'hefb6fa3f0218fef109be0370099f0a2e0aae;
mem[13] = 144'hf779f47bf5a5fa53ff29fe6c06ea01e2056f;
mem[14] = 144'h03d00644047d00f2fb89f7fff65aeb0bf275;
mem[15] = 144'hfcfdffa9062a043407a0030904bdffca007c;
mem[16] = 144'hff1210c419e808970e0f0b2d0d79078a0190;
mem[17] = 144'hf29106620d0ef903fc0006b1fcdafd8f01c6;
mem[18] = 144'h04b00abf01040b890241f0390555f280e8d6;
mem[19] = 144'hff25057cfd2c000f07cb0781fde8060f051d;
mem[20] = 144'h02b4f5cbf37403ecf885f3ddf384f0a2efc4;
mem[21] = 144'h096503f0f88106e80a49020202ad016500f9;
mem[22] = 144'h0f4af28ff0420f9ee67cfa9d1255efbe0507;
mem[23] = 144'h0bd9ff57f48b0b55ff15f31c0c28058df42d;
mem[24] = 144'h0332fd24fbd60133fbe1fbe90415fce7ffe6;
mem[25] = 144'hf8f0017cfdbbf9b5017efbba00f8fca9f987;
mem[26] = 144'hee32fa770594fa14031901bffcfd0795fe38;
mem[27] = 144'hfc75f957f63102c40710056d0267037409df;
mem[28] = 144'h067e0c9e0c7508eb0481fb2c05eeffd9f3bb;
mem[29] = 144'hfce2028603cffbf200cf0590077f06e9ff13;
mem[30] = 144'hede2f7c104d1fb940693105d02ea0e8b0d4c;
mem[31] = 144'hf958f55dfb4efbea007e044c08bd07b209b6;
mem[32] = 144'h0959fcf8fa1b0bc6f6c5f6af00d6f5bbf243;
mem[33] = 144'hff67075b0181fed1022102f5ff62ff4bf5d2;
mem[34] = 144'h05cc0421f8690842ffeaf7a70075fa4dea7a;
mem[35] = 144'h06180160069906a90775092affb000b204a4;
mem[36] = 144'hf9a604ef02c307a6061e00ec034a09ffffbe;
mem[37] = 144'hfca7fa10f7c101b404db004bfe83048f0905;
mem[38] = 144'h03caf931f5270288fda8f1c0fb97f4d9efad;
mem[39] = 144'h069d077dfb76fef20bc002e3fd15017b02b5;
mem[40] = 144'h03a4073e00ea0db8061af5bd0a17faf0f363;
mem[41] = 144'h0161ffd7004609a600bd00aa0918095004a9;
mem[42] = 144'h04ae01f6fb0e0391fdf9f17401f9efcdef63;
mem[43] = 144'hfbf704b6fe5e07ed099c05060657053600bf;
mem[44] = 144'h09c9ee08f506ff40ed8001bdff33f906fe0c;
mem[45] = 144'h077a000ff6e2ff68f8acf63c02e3fc2cfad6;
mem[46] = 144'hf1530c6815d6fc9b0da9196509d914c70f4f;
mem[47] = 144'hf76df6430cb0f2b6f8720b34fb5afd1608e5;
mem[48] = 144'h1222f0d3f31c10c6eef2f5a510aafaf3f6e0;
mem[49] = 144'h0b750109f60d0a3f05e3f3770229fdbcf617;
mem[50] = 144'hfdee0481fae4ff83fd99038efe55fefbfdd9;
mem[51] = 144'hfc96fdcd020e00e40424fa850108fc3bfdfd;
mem[52] = 144'hec6e043a1266f30209f211abff0b15c80d6b;
mem[53] = 144'hfd6cfed30385f6c2fd6c0632f983ff670595;
mem[54] = 144'hfd86ff19fae1fc14016cfede01f5fe71fd49;
mem[55] = 144'hfb4d03d5fc060018fd140031fd7ffacb0083;
mem[56] = 144'h078e02cc000deb1fee0df06ee2c4ee4df517;
mem[57] = 144'h0a45099a0c92fd5e002efd41edecf0a4f50d;
mem[58] = 144'h1106fe8bfa8b0328f2f5f3afe540ebfaf652;
mem[59] = 144'h069007a80ad0056804ee02a1f948f39bfdd6;
mem[60] = 144'h04c0054b099204690d00ff890273002ff7ac;
mem[61] = 144'hf4bf02dbfc16fc5403620659087808be0205;
mem[62] = 144'h01530417f64301e2fea2f65effbbf65bf23e;
mem[63] = 144'h0361037605d0053a05b2fe4c01cb06f00681;
mem[64] = 144'h0a3906ea03480c4f0443f812fa71f2eff116;
mem[65] = 144'hfdfe02ca00760758053802c0035a08780471;
mem[66] = 144'h099f01fe04f1f924f436094b06f2fb3106c1;
mem[67] = 144'hfd6df48dfe1bfa4b0766f4e9ff6bfbb4f7cd;
mem[68] = 144'h050d018afda60097fa7409a0f7c5fb360310;
mem[69] = 144'h0b0ffb4e0369fdc8ff6b067efbc9089ffae8;
mem[70] = 144'hf94d064406c7086a089df2ee017bfa74faa3;
mem[71] = 144'h047907090354f81efb4705d502aa081406c0;
mem[72] = 144'hf1990235f98e026cf833f5f203e3088c0929;
mem[73] = 144'h08e2042e012bff4d076f06b1f91ff553f81f;
mem[74] = 144'h00a9fa2bfd7705d7f91706fbfcf80514ff38;
mem[75] = 144'h02890750ff49f921072f0832fdfdf872fe56;
end

always @ (posedge clk) begin
	q_a <= mem[addr_a];
end

always @ (posedge clk) begin
	q_b <= mem[addr_b];
end

endmodule