module generate_problem(
	input[8:0] problem_index,
	output[23:0] problem
);
	always_comb begin
		case(problem_index)
			9'd000:problem = 24'b000000011011000110100010;
			9'd001:problem = 24'b000000011100000110100000;
			9'd002:problem = 24'b000000011101000110100001;
			9'd003:problem = 24'b000000011110000110100001;
			9'd004:problem = 24'b000000011011001010100011;
			9'd005:problem = 24'b000000011101001010100010;
			9'd006:problem = 24'b000000011011001110100100;
			9'd007:problem = 24'b000000011101001110100011;
			9'd008:problem = 24'b000000011011010010100101;
			9'd009:problem = 24'b000000011101010010100100;
			9'd010:problem = 24'b000000011011010110100110;
			9'd011:problem = 24'b000000011101010110100101;
			9'd012:problem = 24'b000000011011011010100111;
			9'd013:problem = 24'b000000011101011010100110;
			9'd014:problem = 24'b000000011011011110101000;
			9'd015:problem = 24'b000000011101011110100111;
			9'd016:problem = 24'b000000011011100010101001;
			9'd017:problem = 24'b000000011101100010101000;
			9'd018:problem = 24'b000000011101100110101001;
			9'd019:problem = 24'b000000101011000110100011;
			9'd020:problem = 24'b000000101100000110100001;
			9'd021:problem = 24'b000000101101000110100010;
			9'd022:problem = 24'b000000101110000110100010;
			9'd023:problem = 24'b000000101011001010100100;
			9'd024:problem = 24'b000000101100001010100000;
			9'd025:problem = 24'b000000101101001010100100;
			9'd026:problem = 24'b000000101110001010100001;
			9'd027:problem = 24'b000000101011001110100101;
			9'd028:problem = 24'b000000101101001110100110;
			9'd029:problem = 24'b000000101011010010100110;
			9'd030:problem = 24'b000000101101010010101000;
			9'd031:problem = 24'b000000101011010110100111;
			9'd032:problem = 24'b000000101011011010101000;
			9'd033:problem = 24'b000000101011011110101001;
			9'd034:problem = 24'b000000111011000110100100;
			9'd035:problem = 24'b000000111100000110100010;
			9'd036:problem = 24'b000000111101000110100011;
			9'd037:problem = 24'b000000111110000110100011;
			9'd038:problem = 24'b000000111011001010100101;
			9'd039:problem = 24'b000000111100001010100001;
			9'd040:problem = 24'b000000111101001010100110;
			9'd041:problem = 24'b000000111011001110100110;
			9'd042:problem = 24'b000000111100001110100000;
			9'd043:problem = 24'b000000111101001110101001;
			9'd044:problem = 24'b000000111110001110100001;
			9'd045:problem = 24'b000000111011010010100111;
			9'd046:problem = 24'b000000111011010110101000;
			9'd047:problem = 24'b000000111011011010101001;
			9'd048:problem = 24'b000001001011000110100101;
			9'd049:problem = 24'b000001001100000110100011;
			9'd050:problem = 24'b000001001101000110100100;
			9'd051:problem = 24'b000001001110000110100100;
			9'd052:problem = 24'b000001001011001010100110;
			9'd053:problem = 24'b000001001100001010100010;
			9'd054:problem = 24'b000001001101001010101000;
			9'd055:problem = 24'b000001001110001010100010;
			9'd056:problem = 24'b000001001011001110100111;
			9'd057:problem = 24'b000001001100001110100001;
			9'd058:problem = 24'b000001001011010010101000;
			9'd059:problem = 24'b000001001100010010100000;
			9'd060:problem = 24'b000001001110010010100001;
			9'd061:problem = 24'b000001001011010110101001;
			9'd062:problem = 24'b000001011011000110100110;
			9'd063:problem = 24'b000001011100000110100100;
			9'd064:problem = 24'b000001011101000110100101;
			9'd065:problem = 24'b000001011110000110100101;
			9'd066:problem = 24'b000001011011001010100111;
			9'd067:problem = 24'b000001011100001010100011;
			9'd068:problem = 24'b000001011011001110101000;
			9'd069:problem = 24'b000001011100001110100010;
			9'd070:problem = 24'b000001011011010010101001;
			9'd071:problem = 24'b000001011100010010100001;
			9'd072:problem = 24'b000001011100010110100000;
			9'd073:problem = 24'b000001011110010110100001;
			9'd074:problem = 24'b000001101011000110100111;
			9'd075:problem = 24'b000001101100000110100101;
			9'd076:problem = 24'b000001101101000110100110;
			9'd077:problem = 24'b000001101110000110100110;
			9'd078:problem = 24'b000001101011001010101000;
			9'd079:problem = 24'b000001101100001010100100;
			9'd080:problem = 24'b000001101110001010100011;
			9'd081:problem = 24'b000001101011001110101001;
			9'd082:problem = 24'b000001101100001110100011;
			9'd083:problem = 24'b000001101110001110100010;
			9'd084:problem = 24'b000001101100010010100010;
			9'd085:problem = 24'b000001101100010110100001;
			9'd086:problem = 24'b000001101100011010100000;
			9'd087:problem = 24'b000001101110011010100001;
			9'd088:problem = 24'b000001111011000110101000;
			9'd089:problem = 24'b000001111100000110100110;
			9'd090:problem = 24'b000001111101000110100111;
			9'd091:problem = 24'b000001111110000110100111;
			9'd092:problem = 24'b000001111011001010101001;
			9'd093:problem = 24'b000001111100001010100101;
			9'd094:problem = 24'b000001111100001110100100;
			9'd095:problem = 24'b000001111100010010100011;
			9'd096:problem = 24'b000001111100010110100010;
			9'd097:problem = 24'b000001111100011010100001;
			9'd098:problem = 24'b000001111100011110100000;
			9'd099:problem = 24'b000001111110011110100001;
			9'd100:problem = 24'b000010001011000110101001;
			9'd101:problem = 24'b000010001100000110100111;
			9'd102:problem = 24'b000010001101000110101000;
			9'd103:problem = 24'b000010001110000110101000;
			9'd104:problem = 24'b000010001100001010100110;
			9'd105:problem = 24'b000010001110001010100100;
			9'd106:problem = 24'b000010001100001110100101;
			9'd107:problem = 24'b000010001100010010100100;
			9'd108:problem = 24'b000010001110010010100010;
			9'd109:problem = 24'b000010001100010110100011;
			9'd110:problem = 24'b000010001100011010100010;
			9'd111:problem = 24'b000010001100011110100001;
			9'd112:problem = 24'b000010001100100010100000;
			9'd113:problem = 24'b000010001110100010100001;
			9'd114:problem = 24'b000010011100000110101000;
			9'd115:problem = 24'b000010011101000110101001;
			9'd116:problem = 24'b000010011110000110101001;
			9'd117:problem = 24'b000010011100001010100111;
			9'd118:problem = 24'b000010011100001110100110;
			9'd119:problem = 24'b000010011110001110100011;
			9'd120:problem = 24'b000010011100010010100101;
			9'd121:problem = 24'b000010011100010110100100;
			9'd122:problem = 24'b000010011100011010100011;
			9'd123:problem = 24'b000010011100011110100010;
			9'd124:problem = 24'b000010011100100010100001;
			9'd125:problem = 24'b000010011100100110100000;
			9'd126:problem = 24'b000010011110100110100001;
			9'd127:problem = 24'b000100001100000110101001;
			9'd128:problem = 24'b000100001100001010101000;
			9'd129:problem = 24'b000100001110001010100101;
			9'd130:problem = 24'b000100001100001110100111;
			9'd131:problem = 24'b000100001100010010100110;
			9'd132:problem = 24'b000100001100010110100101;
			9'd133:problem = 24'b000100001110010110100010;
			9'd134:problem = 24'b000100001100011010100100;
			9'd135:problem = 24'b000100001100011110100011;
			9'd136:problem = 24'b000100001100100010100010;
			9'd137:problem = 24'b000100001100100110100001;
			9'd138:problem = 24'b000100011100001010101001;
			9'd139:problem = 24'b000100011100001110101000;
			9'd140:problem = 24'b000100011100010010100111;
			9'd141:problem = 24'b000100011100010110100110;
			9'd142:problem = 24'b000100011100011010100101;
			9'd143:problem = 24'b000100011100011110100100;
			9'd144:problem = 24'b000100011100100010100011;
			9'd145:problem = 24'b000100011100100110100010;
			9'd146:problem = 24'b000100101110001010100110;
			9'd147:problem = 24'b000100101100001110101001;
			9'd148:problem = 24'b000100101110001110100100;
			9'd149:problem = 24'b000100101100010010101000;
			9'd150:problem = 24'b000100101110010010100011;
			9'd151:problem = 24'b000100101100010110100111;
			9'd152:problem = 24'b000100101100011010100110;
			9'd153:problem = 24'b000100101110011010100010;
			9'd154:problem = 24'b000100101100011110100101;
			9'd155:problem = 24'b000100101100100010100100;
			9'd156:problem = 24'b000100101100100110100011;
			9'd157:problem = 24'b000100111100010010101001;
			9'd158:problem = 24'b000100111100010110101000;
			9'd159:problem = 24'b000100111100011010100111;
			9'd160:problem = 24'b000100111100011110100110;
			9'd161:problem = 24'b000100111100100010100101;
			9'd162:problem = 24'b000100111100100110100100;
			9'd163:problem = 24'b000101001110001010100111;
			9'd164:problem = 24'b000101001100010110101001;
			9'd165:problem = 24'b000101001100011010101000;
			9'd166:problem = 24'b000101001100011110100111;
			9'd167:problem = 24'b000101001110011110100010;
			9'd168:problem = 24'b000101001100100010100110;
			9'd169:problem = 24'b000101001100100110100101;
			9'd170:problem = 24'b000101011110001110100101;
			9'd171:problem = 24'b000101011110010110100011;
			9'd172:problem = 24'b000101011100011010101001;
			9'd173:problem = 24'b000101011100011110101000;
			9'd174:problem = 24'b000101011100100010100111;
			9'd175:problem = 24'b000101011100100110100110;
			9'd176:problem = 24'b000101101110001010101000;
			9'd177:problem = 24'b000101101110010010100100;
			9'd178:problem = 24'b000101101100011110101001;
			9'd179:problem = 24'b000101101100100010101000;
			9'd180:problem = 24'b000101101110100010100010;
			9'd181:problem = 24'b000101101100100110100111;
			9'd182:problem = 24'b000101111100100010101001;
			9'd183:problem = 24'b000101111100100110101000;
			9'd184:problem = 24'b000110001110001010101001;
			9'd185:problem = 24'b000110001110001110100110;
			9'd186:problem = 24'b000110001110011010100011;
			9'd187:problem = 24'b000110001100100110101001;
			9'd188:problem = 24'b000110001110100110100010;
			9'd189:problem = 24'b001000001110010010100101;
			9'd190:problem = 24'b001000001110010110100100;
			9'd191:problem = 24'b001000011110001110100111;
			9'd192:problem = 24'b001000011110011110100011;
			9'd193:problem = 24'b001001001110001110101000;
			9'd194:problem = 24'b001001001110010010100110;
			9'd195:problem = 24'b001001001110011010100100;
			9'd196:problem = 24'b001001001110100010100011;
			9'd197:problem = 24'b001001011110010110100101;
			9'd198:problem = 24'b001001111110001110101001;
			9'd199:problem = 24'b001001111110100110100011;
			9'd200:problem = 24'b001010001110010010100111;
			9'd201:problem = 24'b001010001110011110100100;
			9'd202:problem = 24'b001100001110010110100110;
			9'd203:problem = 24'b001100001110011010100101;
			9'd204:problem = 24'b001100101110010010101000;
			9'd205:problem = 24'b001100101110100010100100;
			9'd206:problem = 24'b001101011110010110100111;
			9'd207:problem = 24'b001101011110011110100101;
			9'd208:problem = 24'b001101101110010010101001;
			9'd209:problem = 24'b001101101110011010100110;
			9'd210:problem = 24'b001101101110100110100100;
			9'd211:problem = 24'b010000001110010110101000;
			9'd212:problem = 24'b010000001110100010100101;
			9'd213:problem = 24'b010000101110011010100111;
			9'd214:problem = 24'b010000101110011110100110;
			9'd215:problem = 24'b010001011110010110101001;
			9'd216:problem = 24'b010001011110100110100101;
			9'd217:problem = 24'b010010001110011010101000;
			9'd218:problem = 24'b010010001110100010100110;
			9'd219:problem = 24'b010010011110011110100111;
			9'd220:problem = 24'b010101001110011010101001;
			9'd221:problem = 24'b010101001110100110100110;
			9'd222:problem = 24'b010101101110011110101000;
			9'd223:problem = 24'b010101101110100010100111;
			9'd224:problem = 24'b011000111110011110101001;
			9'd225:problem = 24'b011000111110100110100111;
			9'd226:problem = 24'b011001001110100010101000;
			9'd227:problem = 24'b011100101110100010101001;
			9'd228:problem = 24'b011100101110100110101000;
			default:problem = 24'b0;
		endcase
	end
endmodule
