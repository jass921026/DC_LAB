`timescale 1ns/1ns

module wt_fc1_mem0 #(parameter ADDR_WIDTH = 11, DATA_WIDTH = 144, DEPTH = 1024) (
input wire clk,
input wire [ADDR_WIDTH-1:0] addr_a, 
input wire [ADDR_WIDTH-1:0] addr_b, 
output reg [DATA_WIDTH-1:0] q_a,
output reg [DATA_WIDTH-1:0] q_b
);

reg [DATA_WIDTH-1:0] mem [0:DEPTH-1];

initial begin
mem[0] = 144'hfff600c10149020b0157fd370041fbd5fda2;
mem[1] = 144'h021201b0029e02b50278fd0cff6ffc50fdad;
mem[2] = 144'hfe70fe04ffac0197fe77f5950200fddefed2;
mem[3] = 144'h024f013301ca02afff42fcc402a40052ff92;
mem[4] = 144'h013aff95018900e30004fd1801ae01c6fd67;
mem[5] = 144'h008cfabdfb5402a9012501befc81f564eff5;
mem[6] = 144'h011effe8ff560159ff29fe6102ebffdb007e;
mem[7] = 144'hfe12fddcfd5cfe8afc86fb19027b015a001e;
mem[8] = 144'hfec2ff67000a0190017afe18ffd2fdf50013;
mem[9] = 144'h00ebfdc5013f011800d0fde101640058fedc;
mem[10] = 144'h002dff31ff8a01b000f8fc99004efefefd11;
mem[11] = 144'hffbdfda0fef400bff9a6014e0058fb10fbc2;
mem[12] = 144'h0072015a02ce0171ffb6fe54ffc0004efd7a;
mem[13] = 144'hfea3fe63004afe890101ffcaffd201bafe49;
mem[14] = 144'hfee508ad07fc01e9fd27ff00041401b001b9;
mem[15] = 144'hffdb01de025a036a015efb9001b8fdb1fe8b;
mem[16] = 144'h01360039ff39feb8fe89018c0036feb0ffd5;
mem[17] = 144'h0145017a0017fff400d7ff6d005f00b90083;
mem[18] = 144'hfe1100240039ff080151015800afff50fff4;
mem[19] = 144'hffc0008eff910106ff52016e0066fea60054;
mem[20] = 144'hfe4f00f90006ff38ffcd01310170fdd4fe9a;
mem[21] = 144'h007bff660126001ffe62ff02ffc00064ffa8;
mem[22] = 144'hff97fdc50026006ffe0cff5f003bff43001e;
mem[23] = 144'hfdeaff5fffb20107fdd800e4fee7ffdc00c1;
mem[24] = 144'hfe6f00f0fdbc010c00c6014afdceffd6000a;
mem[25] = 144'h0061ff87011affa1ff1ffec700c0ffe9fe45;
mem[26] = 144'h0189ff92ff410024ffaa011efdc6ff8dffbd;
mem[27] = 144'h0049feea0041003d00f0ff75fe84fee8fec7;
mem[28] = 144'hffdf000700fb01db004a01680091ff670022;
mem[29] = 144'h00b2fe5ffe89fea8006d0005fff8ff470112;
mem[30] = 144'h005dff43009000e6fe52004001060145fee3;
mem[31] = 144'hfe76fe3f0061012b002bfff6ffd9fe3200ce;
mem[32] = 144'h0050ff30fe64013400dcfe99ffb00189ffb5;
mem[33] = 144'hfeb80104feabff9c005100deff2efe700162;
mem[34] = 144'hfeeffff60042ff11006701d90159fe51ff56;
mem[35] = 144'hfec6ffeaff8dfdc70070ff87fe5a0152ff0b;
mem[36] = 144'hff2a013a0046ffc701830026fef5ff34fff5;
mem[37] = 144'hff98fde20089015cff94fdf3ffe2fe6bff92;
mem[38] = 144'h016c005afec10000004bff55feb501a7ff5c;
mem[39] = 144'hff95ff78fef10049ff89fe66002e00040178;
mem[40] = 144'h00220088febe0149fee6006cfdcdfee2fecd;
mem[41] = 144'hff08ff9100f3012d00ff00a401d6fe6b0020;
mem[42] = 144'h014900d1ff7dff77ffae01980037002f00ac;
mem[43] = 144'hfe8a0120008bff9b011bfe7201bbff56ff6a;
mem[44] = 144'hfffa0053ffd2fef400fe016a00b1ff58ff4a;
mem[45] = 144'hff0200da01180047019dffd0fed900be0081;
mem[46] = 144'h00f10049fdd40096ff70015dff8700e000b3;
mem[47] = 144'hff9d0094febe00d3ffef00c5fe90009affd8;
mem[48] = 144'h009fffaf003aff50fe3e003900bbfea70095;
mem[49] = 144'hfea3000200be00fbfedbff35fe13ffdffe97;
mem[50] = 144'h001cfec7ff9b0095fea9fd80fd78ff3b0032;
mem[51] = 144'h007fff19fdf7fe13ff1afe60fec50033fed1;
mem[52] = 144'hfef2fe68fda7fd7bfe67ff1eff5bff8700d2;
mem[53] = 144'hfe92fe65ff1c00fc004e00d5ffa4fe2cfe1c;
mem[54] = 144'hfde0fd81004fff63fd7700fefe12009dff8b;
mem[55] = 144'h0002ffa1fff1fe7cff24feb3ffbbfe760088;
mem[56] = 144'hfdaffe54003afdbd00a7ff53fe2500ecfef5;
mem[57] = 144'hfe21007dfe0eff7effbbfe4600f4007aff9b;
mem[58] = 144'h002cfe79fe74ff10ff7cffdafdf3006efd7c;
mem[59] = 144'hfdf4fe06ffa6ff4bfd7d010c0077ff8aff23;
mem[60] = 144'h018dfeeffe9b0068002fff4600c1003ffe31;
mem[61] = 144'h00310156ffd00089ff450097fe58febb01a5;
mem[62] = 144'hfd7200feffc3ffc3fdd200fbffa7ffa10020;
mem[63] = 144'hfdb3fe73fde2ff93ff65fffbfe88fdc6ff21;
mem[64] = 144'hff71fd37fe80ffd3fe14fb7efddc017fffd8;
mem[65] = 144'hfee6fe6aff150003fffffec3fed4ff460258;
mem[66] = 144'hfb10ffe20018ff1ffe900716007d02030005;
mem[67] = 144'hfe21fcc6febc017a00bfffd0fe8bfe280235;
mem[68] = 144'hfe3bffdafe4a026d00daffaeff97ff160200;
mem[69] = 144'hfedbffdffc4efe770257fd7902b700b90506;
mem[70] = 144'hfe0efe8d0286027301beff87fffc027702c0;
mem[71] = 144'hff1bff52019b04fc03e602ba01c703bdff7b;
mem[72] = 144'hfe42ffcb007c0116fe4200a7feb2016100d1;
mem[73] = 144'hfdc5ff96ff96fe6dff86fd62fd1ffeb00207;
mem[74] = 144'hfd34ffee0002ff0b0198ffbefdd4ff8a0192;
mem[75] = 144'hff44fe0affc60120fca801a3002bffc90403;
mem[76] = 144'h004d0157feb3feecffe4ff6200ef014b0058;
mem[77] = 144'h000fff0eff70fe98fe6f014dff4a00d60039;
mem[78] = 144'hfeeffd45fb7cfd61f897fb21fd53fd1bfe2e;
mem[79] = 144'hff48fbcaff200174ff6efea8fdb4028a017b;
mem[80] = 144'hff07fddbfeccfff1005efff4fe3600740104;
mem[81] = 144'h00e50045ff8f008e00f0014fff25fefcfe82;
mem[82] = 144'h016cfecb000cff74fe4e0120ff97ff1dff89;
mem[83] = 144'hfdbdfe810019fef6fddcffe5fe6d00d4fe98;
mem[84] = 144'hfe79ff23fde600470043fedefdbeff69fe33;
mem[85] = 144'hff5100400162fe72fea000780149ff27fe92;
mem[86] = 144'hfdccfe50fe8500d6fe04010ffef4fe1d006e;
mem[87] = 144'hfe73009b0180017f0096ffc0fe0b0225fe8c;
mem[88] = 144'hfe370111fdc9ff74ff96ffa6ff33fe4b014d;
mem[89] = 144'h017afe76fe5600d3001e01c90151fe8effee;
mem[90] = 144'h01720151ff3bfe5500b4013100cdffd0006c;
mem[91] = 144'hfddd0075ff95ff77ff9e00ccfe0cff9afe69;
mem[92] = 144'h001c014afe840148fffe0115005300590175;
mem[93] = 144'h014e00cb0106ff03ff78fe5f01afff62ff98;
mem[94] = 144'hff23ff6c0131fde60101005a008cfdceffdc;
mem[95] = 144'h014f009d011efe88ffb3fe6dfe61ff75fe10;
mem[96] = 144'hfc3001c3047402f30245037cfbe90158fec5;
mem[97] = 144'hfd4900cf039b03c002e20405fc0dff510001;
mem[98] = 144'hfc8e004a01f003140192035201a301fb0335;
mem[99] = 144'hff39012301c4021704200392001100f3fec0;
mem[100] = 144'hffd90185014b034a01080315fdd400db0033;
mem[101] = 144'h00b902000023fda30198fffa00b307e009b1;
mem[102] = 144'h00430179010302d50237013601bc0121fda0;
mem[103] = 144'hffcaff26fe7f000dff6b014b025e00e10034;
mem[104] = 144'hfd2f01ae0412051503af02beffb7013cfde2;
mem[105] = 144'hfe69021c0448033002190374fcf7fd12fe32;
mem[106] = 144'hfc02fecb02c90435040a031cffc7ff14ffbb;
mem[107] = 144'h00e9016803bbfe87fd51fd47008702b1031f;
mem[108] = 144'hffb100b500a5011d007e004afeb7024a020c;
mem[109] = 144'h00cf01260016ff5fff70ffbc00870122ffc7;
mem[110] = 144'hfd86fcdbffd2051c02de039cfbd6ffb40188;
mem[111] = 144'hfbfb025003e5035201c80419fe0000ebffa8;
mem[112] = 144'hffcbfebe001f012f00edff66ff96fe5affcb;
mem[113] = 144'hfee7ffd5fe4effabfedcfe45ff17ff06fe82;
mem[114] = 144'h0080fe9d006600b0fe5900e2023bffab0144;
mem[115] = 144'hff1afe510039006e002dfeb70177ff1eff61;
mem[116] = 144'hfef3ffe0003f0176013bff63009400b5009c;
mem[117] = 144'h00190127fdc40000fefdfed9005301770108;
mem[118] = 144'h0011fe14012eff1eff8dffadfde9fee80076;
mem[119] = 144'hfffcfe29ffbbfef9007aff2fff0400b6014a;
mem[120] = 144'h0050fe00010700defdd9fe1fffd5ffcdfe77;
mem[121] = 144'hff50015dfee3fec6006aff90010101b7fe89;
mem[122] = 144'hff03015cfebc005bfdd8fe2201f4023cffa6;
mem[123] = 144'hff7200c1ff52fedfffc0fea2014800b6fdec;
mem[124] = 144'hfe800197ff5b018c019e017aff4eff5f0038;
mem[125] = 144'hff8600d200e8fe8e0171feaefeaf005d015d;
mem[126] = 144'h0077002f0164fe35fee200c0fdf500f2fe1f;
mem[127] = 144'hfff4005500e90114fef2ff99006bfdefffbf;
mem[128] = 144'h01be012afc8bff4500e102d8021a03eaff7a;
mem[129] = 144'h027dff9efce1fe2c00e703de03fc036a00f9;
mem[130] = 144'h041b003cfd400049039409a70208fed2feba;
mem[131] = 144'h01dc0252014afe72fee2012b018a0239fee2;
mem[132] = 144'h03100203000f0013ffc10135021702caff97;
mem[133] = 144'hfed103090510fd42fe44ffbaff0103ec0ade;
mem[134] = 144'h02160104004b0072025e021e025b0046ffdd;
mem[135] = 144'h029a0175011f01a5009d02190060fd41006a;
mem[136] = 144'h0234fff00094ff960233013f01730329ffb1;
mem[137] = 144'h02aa007bff09ff0affc1016500ae03f20264;
mem[138] = 144'h016d03fe01bdfde8fdb8012600f5007b0045;
mem[139] = 144'h001aff9afd2d048c0711013d0146001f009e;
mem[140] = 144'hffa6ff11000000d2003f00faff0bfe83ff9b;
mem[141] = 144'hff1800e0fe72ffdd00cbfe6fff8cfefcfea6;
mem[142] = 144'h0207ffd2fe65fe3600c7003901a60195ff30;
mem[143] = 144'h010103080071fdf501a1017702d503f50100;
mem[144] = 144'h04b1016202880089fd5af76802c0ffe702d6;
mem[145] = 144'h018001c8050c02edfea3fcc6033d00e00532;
mem[146] = 144'h017b0394027afe6efe13f96f0213fc6efd61;
mem[147] = 144'h003702a00235028affb2ff32047802240357;
mem[148] = 144'h005f014104fb01ed00a7fea802d1011600ea;
mem[149] = 144'h0034fd0bfd5d01a60244009dfdf9f5e1f02c;
mem[150] = 144'h0377028f035b00e30137ff680301fe3103e0;
mem[151] = 144'h01d702ee015b038b013602090115ff07ff33;
mem[152] = 144'h000d0080048effc9ff60fe030240023303da;
mem[153] = 144'h029202be0299030afde1f9f901c8017900a1;
mem[154] = 144'h02ed0480024e026400bffd87024402e60284;
mem[155] = 144'h00ae014afcb5f849f812021bff61fb99f954;
mem[156] = 144'hffa7028702e90010012c00ab0147fd49fcd6;
mem[157] = 144'hff9e019bfe3301440117fec7ff59009ffe3c;
mem[158] = 144'hffdb023c01f9003ff9acfa9903c805e30479;
mem[159] = 144'h00910470032d00eaff96fc03019400a301e4;
mem[160] = 144'hfce6fea5fc59ff42fe390049fc9402890051;
mem[161] = 144'hfefffe4fff3ffe570011fefdfd0cfff703b5;
mem[162] = 144'hfbfe004affa5023e007d044bffe001420174;
mem[163] = 144'hfd760040ffe0fe2bfe100004fecd01040277;
mem[164] = 144'h00b901400139001eff8f0184fd8e023f025c;
mem[165] = 144'h01c401e90113fca3027cff6b03e103ab0553;
mem[166] = 144'h0025009101580173006800e1fd1e021f02af;
mem[167] = 144'h000e012e01ca031400fb038aff89001802fd;
mem[168] = 144'hfda0009dfc79fdc4014c00eafc1400ed017a;
mem[169] = 144'hfd95ffa9ff7cfdacfe16ff2dfba601da0315;
mem[170] = 144'hff37ff57ffabfdb200dc0062fbf200e80304;
mem[171] = 144'h003d019afe26fe9cfe5a0168002703b6039c;
mem[172] = 144'h00adfeaffeec001100fa00bafe000098fffc;
mem[173] = 144'hffe8ff5201ab0009feccff0d00ea007a01ab;
mem[174] = 144'h01b5fd8efba1fece01caffa3fb39006901db;
mem[175] = 144'hfe460139fead0091fe0100bffc3b009501ec;
mem[176] = 144'hfe9efe86fdf6ffcefe77ffdffffe001aff53;
mem[177] = 144'hff0c0049ff58feb6ff61fe9dfe1dfebf00a2;
mem[178] = 144'h013601ccfdc2fdc1ffcb002901720102010b;
mem[179] = 144'h016c00500166ff98fe92fe4dff5f0161fee2;
mem[180] = 144'hff4dfefdfffaffe4fe770017fe1dfddb0159;
mem[181] = 144'h00eaffc9feeb00bffe1cfde80091fde2fffa;
mem[182] = 144'h009c00daffdefedffdc1ffaefe24ff3cff87;
mem[183] = 144'hfe53fdf300a600b40003ff990071ff880144;
mem[184] = 144'h0034009dff2bff9b0073fe2dfe3ffde7ff51;
mem[185] = 144'h0043fed0ff3300d1ff7bff2200fcff95fee0;
mem[186] = 144'hff73ffa9fe260003fe2e000a002101930152;
mem[187] = 144'hffd101b000e900c80068fed80220010efe00;
mem[188] = 144'h015fffeb00d9ff1f0032fe2200edfe550126;
mem[189] = 144'h004cfe42ffbc007600b0ff7d009f00b500bd;
mem[190] = 144'hffdeff8dffaeff180117009fff13febf012b;
mem[191] = 144'h00b7ff0bfdf0011e01010146fe950123fe18;
mem[192] = 144'h01f50057fe25fea6044f0312027d02f2fde5;
mem[193] = 144'h0080ff4500c8012f0250043e024800f6003f;
mem[194] = 144'h04440203fd64ff2e02e20451005500a4fe27;
mem[195] = 144'h014701d60197fea50108011501de00edfdac;
mem[196] = 144'h01290174fe9c01120231039d023dfff7fe89;
mem[197] = 144'hfe1cff8bff3c021001ed007bfd4c023d0835;
mem[198] = 144'h01a30251fd47ff44011501a0013f0262fe7a;
mem[199] = 144'h029400cbfeacfe1efe63ffc6fe00ff5afbd7;
mem[200] = 144'h0123001200e5021601240283038b0024fe3e;
mem[201] = 144'h018b02ec008b00b301ec019701a602db022f;
mem[202] = 144'h026100c600320016008803b001470110fea8;
mem[203] = 144'h0146fd82011804e80276fde800f901000066;
mem[204] = 144'hfe8afea0fee7ff6eff61016aff5000defee3;
mem[205] = 144'h00820161ffb8ff560029fe9c0073006c01df;
mem[206] = 144'hfda2fea2005d0150009701df0397ffadfede;
mem[207] = 144'h002c00c8ffbcfe6bffda0154014dff9cff6e;
mem[208] = 144'h01b8ff43ff6dfddcfbddfde302b1009c008c;
mem[209] = 144'h0334fe22fcd8fc9efde0ffc30163005902d9;
mem[210] = 144'h00a3fe0bffc4fd2800ea0268fefe00de0009;
mem[211] = 144'h00f30003ff9cfdfffd5301e7017bfeab0022;
mem[212] = 144'h0282004d0167fe7ffe3400f501e701c1029a;
mem[213] = 144'h002d021b03ef0328fde202bd0282019c0436;
mem[214] = 144'h010602b50210fe41ffe40271020601e70221;
mem[215] = 144'h0090020f01c402c903d2025b012e00e2feaf;
mem[216] = 144'h02fbfccdfda4fdf1006300db02c3013b005a;
mem[217] = 144'h02e8fee5fdb3fb63fc95fff6020602c50199;
mem[218] = 144'h010dffd4009dfed3fcab0141ffc7005f0445;
mem[219] = 144'hfe80fd770021025c078d033600a5023b03fa;
mem[220] = 144'hfea4ff0effbf0180ff3500f2ff75ff7efd87;
mem[221] = 144'hffcafe620084fe58fe7c0157ff85003bfec5;
mem[222] = 144'h0399fd4cfaccf994fc96014503f80220ff47;
mem[223] = 144'h0308fdf0fcb1fe7c0018003a012701d500c7;
mem[224] = 144'hff0802bf050c0407fca2fbd500f4022b03b1;
mem[225] = 144'hff52035b02e302f7febafb77ffe601370475;
mem[226] = 144'h00fc04f70502038efcbbfc9b0214012d01f5;
mem[227] = 144'hfcacff9b038b0199016efe330074028c0589;
mem[228] = 144'hfd8aff6d02ef03d801f8fc72ffa801f30440;
mem[229] = 144'hff7efcb7f711fc6d0079ff8dfe38f64ff0b6;
mem[230] = 144'h006004230571059000d8fddeff8902a100eb;
mem[231] = 144'h01d601480481048003c70178027200e3fe39;
mem[232] = 144'hfd300241036c00dc00eefc85ff300434048d;
mem[233] = 144'hfc85024a014b02c6fdecfd05016001b900f1;
mem[234] = 144'hfd7001b603bf042c00f1fd2f00a903c70456;
mem[235] = 144'h01de02effcfbf80af33000e1010e0001fa15;
mem[236] = 144'hfe7802ab01affef7fefe01b0ff02fea601fb;
mem[237] = 144'hfff900ea00ae013000d7fe9dff53000c00bc;
mem[238] = 144'hff5700e604500296fddefaf4ff3f0453058a;
mem[239] = 144'hff1f03b6043b0227feaafe3200ee033b0481;
mem[240] = 144'hfd6dfdfeffce0163039c0298fdb5008afd4b;
mem[241] = 144'hffd1fdbeffa00245020e0251fd4efcca0006;
mem[242] = 144'hfabbfedd02b2040403e60572fea100800627;
mem[243] = 144'hfdb8fd69fef1001a033402c6fcd7fd550130;
mem[244] = 144'hffecff3dff5f024303340356ffe7fee40147;
mem[245] = 144'h026105ba0301014e0155009907370c560cb3;
mem[246] = 144'hfd60003700b601bd0171ffd70061fe9b008b;
mem[247] = 144'h00bc0065ff26018400d30109ffe401f20321;
mem[248] = 144'hff32004efe4800b5019e02ddfc840089fe70;
mem[249] = 144'hfde4fd160054003b02dd044bfc69fca4fd74;
mem[250] = 144'hfd3cfdacfdc8008700ee012dfd04fdc8ffbb;
mem[251] = 144'hffed0354038e06bf06c000cafff0046d0de1;
mem[252] = 144'h0012fe43fdb7fe9201b4ff730128008d0193;
mem[253] = 144'hff8401b6ff300037fef1012f0055fec0016c;
mem[254] = 144'h01f1fc89fae400ae04a7034ffbcbf97dff60;
mem[255] = 144'hfdceff5cfe7c02f20068015aff190071ff8b;
mem[256] = 144'h008e01d900d500b1020505a000290191ffad;
mem[257] = 144'h018503d3fff803ab04be0475030700ff000c;
mem[258] = 144'h03b2ff4d02160172018d03b00235fedf0280;
mem[259] = 144'h0169006cff2f03970167001a02f700a6011e;
mem[260] = 144'hff6afef2fefa01d1015c017801790154fe5f;
mem[261] = 144'hffd40035ff71ff920196ff6301bb00f20049;
mem[262] = 144'h00e300dcff68fdfeff9400a3016dfd4cfca4;
mem[263] = 144'hffdb00a3fda000b3fce1ff4000f2fed4ffbd;
mem[264] = 144'h01b7023aff6003ff044201ab02b3ffff01f0;
mem[265] = 144'h0274025a000b020f02c8033f020cfe87fdff;
mem[266] = 144'h01dd008cff9102870157ffd3034a025bfdff;
mem[267] = 144'h0246027a019800fdffacffa600b70053fe9a;
mem[268] = 144'h01b7ff68ff26ffceff7eff4600d6ffe8fecd;
mem[269] = 144'h004bfeb5ffddff7bfeaa01bbff4afe6801a7;
mem[270] = 144'hff59017c011603f0089b069dff70ffef0120;
mem[271] = 144'h025803c20147022703bd004102c000bd022e;
mem[272] = 144'hfafdff80020501ca046f0141fb980232ffdb;
mem[273] = 144'hfe3e01580246013803a500c2fde3002aff1f;
mem[274] = 144'hfc0b025f00fc042afecefe0e005b01ff02e9;
mem[275] = 144'hfbdeff5002e000c6010bff39fbe0ff7f022d;
mem[276] = 144'hfd0e0098feb4038e020afdc7fdc6027e027b;
mem[277] = 144'h030300fdffdbfc9d002ffec80453032c01b2;
mem[278] = 144'h000d004c00be0038002bfcdd01d00169fdba;
mem[279] = 144'hfeb2fe98fffd016c011ffeae027b038602d1;
mem[280] = 144'hfec9ff1000080102016d016bfdfbff5401ba;
mem[281] = 144'hfeb10047fe95036802bbfe05fc93fecffd84;
mem[282] = 144'hfe41ff9dfe2802e8025c0001fdf4ff20000a;
mem[283] = 144'h01ec0219fff301c9f946fd3602890479fe09;
mem[284] = 144'hffa800de0010fea8ffa1fe6000e9006c0138;
mem[285] = 144'h01bd0083006eff21002fffcaff1efff00100;
mem[286] = 144'hfe2f005dff7e029e07c8032bf935fce40005;
mem[287] = 144'hff0b01bc02a0030903e9013cfc7300e401f7;
mem[288] = 144'h022afe5300f20354009c01d9febc0064ff74;
mem[289] = 144'h026d004f025b028b025000bfffef01290211;
mem[290] = 144'h008bffbe0320019201150ac100ba0379fec4;
mem[291] = 144'h0089fdd00356011502170197ff19020802aa;
mem[292] = 144'hff96fec80112007a0059021c0038ff6c0083;
mem[293] = 144'h02c301dbfe0ffeaf01c6000204750185059f;
mem[294] = 144'hffa1ffe903af04ad03ba03c8fead0024fdf2;
mem[295] = 144'hfe76025a046e041f018d058e010effdefd3a;
mem[296] = 144'h01f90021003c03190002019cfe14ff000139;
mem[297] = 144'h0042008b002fffcb027a0099fe4300baff39;
mem[298] = 144'h0298fe25021703c300de02a00026ff8601da;
mem[299] = 144'hfebb017003d1fc50fc3401ab01410424011f;
mem[300] = 144'h0167ffffff8701a401ad00be028000740002;
mem[301] = 144'hfe35ff6dff05fe82ff860141fead01d100e4;
mem[302] = 144'hff74fe8efc4600ff0307ffd5ffb9fc5c0239;
mem[303] = 144'h01a6fdc900dcffe9031f0344fe9300360116;
mem[304] = 144'hff52ff6cfe73ffaaffe60045ff120139fe6b;
mem[305] = 144'hffbdfe44012bfe80fe29ffad003cfeabff16;
mem[306] = 144'h0004fffefdb300f5010bfe2ffffffff4ff78;
mem[307] = 144'h007dffb4ffe2fddefe22ff4b00acffbafe6a;
mem[308] = 144'hfecf0172002e0004ff5d0010fef1015cfe14;
mem[309] = 144'hfe720059fff2ffa0fe75fe66fed0016dff55;
mem[310] = 144'h0017fdc400fefe55fed300b5ffb7ff29008e;
mem[311] = 144'hffe5febd00b50158ff2bfe1eff5dff53005a;
mem[312] = 144'h005afe81ff79febefeef00a3ffac014b011d;
mem[313] = 144'hff890176fdd5014e00df015afe74002effcc;
mem[314] = 144'h0093003dffe6fe00ffadfec7fff5ff8efe18;
mem[315] = 144'h012e003001450095002f0069fe0dfe47ffc6;
mem[316] = 144'hff36fe9d007d013dffdd01cf017bfeedffb5;
mem[317] = 144'hfefcffcdff42ff96fe2100f3005aff00ff56;
mem[318] = 144'hff37ff97fe5500c7ff680164ffd0ff7bff11;
mem[319] = 144'hfde600b000320040feb8fdd6fe12011cfe2b;
mem[320] = 144'h0336fb92fdebfda10001fe5f003ffc4efcd9;
mem[321] = 144'h0265ff4ffd16ff20ffef01cb01e4ff50fd75;
mem[322] = 144'h0169fd47fd9c000e00a9fbc1fb9bfd0d0144;
mem[323] = 144'h04fafcedfc4efead007201270156fbea00a1;
mem[324] = 144'h034effab0007fd8a019e0041020bfc5dff9d;
mem[325] = 144'h01cd04b0040e06f00325026401360404048f;
mem[326] = 144'h01d8fe8bfebc01130068ff52002dfe75fe60;
mem[327] = 144'h009dfeba023700340127fc7efde1ff36030e;
mem[328] = 144'h03c6ff0efd73fd53ff200078ffcdfc5dfe0f;
mem[329] = 144'h04c7ff5afeb1fd35019e020e00defe450084;
mem[330] = 144'h0263ff7bff58fec900edfecc012cfed1008d;
mem[331] = 144'hfee7feec03d90981081d00f4fe7afd6808f9;
mem[332] = 144'hfe540055002cfef8ff7900aa01c7ff51fe49;
mem[333] = 144'hfe74feb100d5007200b801440130fec3fee0;
mem[334] = 144'h014001c3feb0f9c0fcc2029f03e9ff7ffb65;
mem[335] = 144'h025fff4afc58ff0e00b7008a0137ff330024;
mem[336] = 144'h0169019cfddffe0f036d074b005300b4ff78;
mem[337] = 144'h0290011efcd5fd05033105aa009c01a201c1;
mem[338] = 144'h00cf01d5ff8efe5704d60989002801c4ff13;
mem[339] = 144'h0134fff3fdd8fff2ffed0204025a006b00bd;
mem[340] = 144'h01be016a00d8fd98ffde0156ffa702bc01db;
mem[341] = 144'h019901a20670ff670061ff95001a076510fb;
mem[342] = 144'h0047016fff580035ffc7054b0142009ffdb0;
mem[343] = 144'h022101bc0171fe37ff0c007c0011fee3ff0e;
mem[344] = 144'hffc60019fed2ffde010e04e4005c016f0033;
mem[345] = 144'h023100c40002feec00ad06c2024c00880071;
mem[346] = 144'h01f80177ffd1ff07fded031a01ac01190299;
mem[347] = 144'hffd3fe8700c408c50a62000f01f0056e037d;
mem[348] = 144'h0086fd83fef8fead0113ff350082fdac0032;
mem[349] = 144'h00a000b4fed4018dff40fe84fe48ffe3010c;
mem[350] = 144'h0242fdccfb2afff306ae051dfe77ff82fc50;
mem[351] = 144'h03590194fdadfea10278064b00cf0250000a;
mem[352] = 144'hffccff7aff25007e018b009cfe44fcb4ff1f;
mem[353] = 144'h00470077fe7bfef40103ffacfc6afdb8fe94;
mem[354] = 144'h004ffe66fdd8fd1d005101bcfc2bfd0cfd6d;
mem[355] = 144'h009b018dffa5fd6efe38ff53fd8afdf5fda9;
mem[356] = 144'h0067ff25fe5ffeb9017901ecffaffd7cfed1;
mem[357] = 144'h0180ffbb00de02c5028900c502ba02d5055d;
mem[358] = 144'h00b10090fe90ffae029b000afc0ffddf0037;
mem[359] = 144'h021afe5dff89fe9c02490053fe6eff9201b6;
mem[360] = 144'hff5e00d0ffb201550073fea8ff0dfe9cfe34;
mem[361] = 144'hff8e01dc014601010271004ffddfffd700a2;
mem[362] = 144'h01e3fe3cfef4fd00ff2301dbfc30fbe7fdd4;
mem[363] = 144'hff97ff22fe700343058600b1fc58ff01ff13;
mem[364] = 144'h014401e6ffbb00ceff15017aff3602ae019f;
mem[365] = 144'hff7500b9ff32ff80ff9afeb6ff4001a2011b;
mem[366] = 144'h00a9fe6b01f20019fd89fc7f001dff1aff22;
mem[367] = 144'hffa1ff7dfd7efd28011901f0fdc6fdb9fc0c;
mem[368] = 144'hfeeafdd500630123ff4b004600c0fe1b007b;
mem[369] = 144'hff92febb014a0118fe72ff61ff82fec6ff52;
mem[370] = 144'h0173fffefebc0160fe3a01b900fd00120008;
mem[371] = 144'h012eff61ffc200790066ff5effad00ee0134;
mem[372] = 144'h00810116015eff480168ff0f017efff4fff9;
mem[373] = 144'hff3bfebdfef400620132feafff4dfe710123;
mem[374] = 144'h012ffedc00aa00140166fe00fec4fe070053;
mem[375] = 144'hff93013dfe1bff12012fff8ffe4cff0f0137;
mem[376] = 144'hfe14001e001affab006cfe4efe6aff2a003d;
mem[377] = 144'hfdf8000c0061fefe00b3016cfe3a01a300c1;
mem[378] = 144'hfe4d009e0096006d002cfee400b5fe63fecd;
mem[379] = 144'hffcbfe0900ac005bffa5fe4c00ff012c014a;
mem[380] = 144'h014a01beff25fe6fff93ff1b01aa0118004b;
mem[381] = 144'h001601b7ffacffd2ff3cff9d001b00000123;
mem[382] = 144'hfef7010bfde0002ffee7ff33fe91fedf00df;
mem[383] = 144'hff5cffd1feb5ff21012b001dfdd0fe45fecc;
mem[384] = 144'hfe97fed0ffd5fee1ff9dff3e00a500f5fd8a;
mem[385] = 144'hfd63fe1e0057ff4c0069fec4ff46005e0038;
mem[386] = 144'hffc0fd320036fe0cfe73ff3dff4a010aff94;
mem[387] = 144'hfd77ff7ffebb001c0032fe99fd9600a9fe85;
mem[388] = 144'hfd7bfce9fdc4ffd6ff5cfe23fd6aff3efee8;
mem[389] = 144'hfe83fef6ff030029ff2efe510126fcc4ff2e;
mem[390] = 144'hfe91fdeeff2e000600c100f100aeffa1feb6;
mem[391] = 144'hfedbfe56ffaffefefefffd99fffb00e9fd99;
mem[392] = 144'hfe79ff51fde3fd11fe5bffaffe79fe1c0029;
mem[393] = 144'hff06ff33ff48fff0002affb9005c01290034;
mem[394] = 144'hfe91fe1dfe51003bfe2400ae0099fdaf00b0;
mem[395] = 144'h005300760089fdecfe02001cfecc0011fddc;
mem[396] = 144'h016f00e4014100aefec5feeafe5c0040ffa3;
mem[397] = 144'h008f0069ff62fe7901ce0163011afff101a9;
mem[398] = 144'hfec7ff65fd50fdc0ff1efeedfcb1fcc1001c;
mem[399] = 144'hfd6cfdeffe81fd66fe19ffaefeb1fedfff63;
mem[400] = 144'h0167fee4fcbffc1efc59fa16fddafe3bfe37;
mem[401] = 144'h021cfcddfdbffe60fe57fc3fffa6ffcb012b;
mem[402] = 144'hfde4fcb1fdc1fd32fc6402eafa15ff9cfe40;
mem[403] = 144'hff9dff75fd82fd1bfcfb0049fed0fd8ffe63;
mem[404] = 144'h019f0116fe46ff24fc61ffdbfe83fe4fff2b;
mem[405] = 144'h0240ffdc02df033f003aff7100e2011e022c;
mem[406] = 144'h0010feb2009dfd65fef5ff35fe95fec60086;
mem[407] = 144'hff77ff9300d500f4021e00d3fde700e201fd;
mem[408] = 144'h00a5fdc3fcb5ff2afed8fe880062fed0febe;
mem[409] = 144'h01af0121feaefb79fbf6ff6effa7ff160382;
mem[410] = 144'hfeacff4afe1cfb6ffddbfc96ff2dff080000;
mem[411] = 144'hfd8efe31fed20008041f0124fca6feecffc6;
mem[412] = 144'h00c1ff6c0081ff03ff760165ff730028ff58;
mem[413] = 144'hffe4007d014a01370000fea8ff2d0141ff15;
mem[414] = 144'h0039fcfafc55fb44fe1bfc1c0219007600d0;
mem[415] = 144'h020dfe39fe76fb79fcc3fd97ffccfe18fdf8;
mem[416] = 144'hfd68ff7bfe780246fe7efd1cfc70fdebffab;
mem[417] = 144'hfc20fd09ff960240ff1efd9bff45005afdf1;
mem[418] = 144'hfc28ff2bffebfde500070081fd71fe57fc0d;
mem[419] = 144'hfd81ff83fe0b017f0032ff45fc36fef5fda9;
mem[420] = 144'hfe1cfc2d017a01abfd5bfe47fc7ffdb1ffb7;
mem[421] = 144'hfd0bfd82fcf4fb73ff1ffedbfe5f007300f2;
mem[422] = 144'hfb64fe4ffe87009bffe1ff7effadfe4afcf2;
mem[423] = 144'hfe31ffeffe0dfe4afd79fda9fe68fe90ff26;
mem[424] = 144'hfd10005dfe76000dfda6fe2bfe2e0004fe98;
mem[425] = 144'hfc3ffee10002017b0140ff61fe36fff5ffc6;
mem[426] = 144'hfc19fdbefddc00d600e4000eff0900f0fca2;
mem[427] = 144'hfc9afe24fd64feedfeedfe15ff23fe57fc7e;
mem[428] = 144'hfe56016300c600e1fe60012dff16ff39ffdc;
mem[429] = 144'h01ba002cff57fea901a2ffedff380188007b;
mem[430] = 144'hffa6ff2b00d90007ff45000bfec1feaa00b2;
mem[431] = 144'hfc89fefafe4e0129ffac007ffcacfea5fd53;
mem[432] = 144'hfe0600ddff12ffe600abfed7fe52ffe10048;
mem[433] = 144'hfff80115ff3f015afdf200e2ff0affcb00b1;
mem[434] = 144'hffacfe9cff65ff80005dff45ff2c0020003e;
mem[435] = 144'hfe0fffafffe0ff450044fe9cffe4ffefff15;
mem[436] = 144'hff59fe72fec4ffbcfe5efefcff43fef2fe98;
mem[437] = 144'h0128fdfd005f0052ffdb00d5ff4200fa01ce;
mem[438] = 144'hfebefe610129ffe0ff98ffddffbdffbfff12;
mem[439] = 144'hffb9feb1fe55feb4ffd0ffc10112011a00e6;
mem[440] = 144'h00c2fe3efeea005700040158fec20144ff2e;
mem[441] = 144'h00ff012efe99ffe1ff4100c0fe41ff23ff8e;
mem[442] = 144'hfdc6fe58fe3afdedff5cfe970015ff2d00ad;
mem[443] = 144'hff83021a003100ae01d1000efeadfee200f0;
mem[444] = 144'h0107fe99fe8b018efe6cfe39009d0105001a;
mem[445] = 144'h00a8ff8800ecfebbfea2fe2d01e1ffd0006d;
mem[446] = 144'hfdda00d8ff6a00a3fdf9fe05007300cf0072;
mem[447] = 144'h0077ffbc00d7ff0efea9ff6bfddaff48fdae;
mem[448] = 144'hff50010fff0efe210059012efdc0ff3aff8f;
mem[449] = 144'hff09fff5ff80febafffeff9dfede0113ff33;
mem[450] = 144'hfeb7005900440119ffbe01aaff7a007ffef1;
mem[451] = 144'h0067fdc5fec0ffdf0108fe9bfde2002ffe5b;
mem[452] = 144'h01770012fde7fe730030fed70038fe37fe84;
mem[453] = 144'h0170ff02ff9a00060037ff0effc3ff53ff39;
mem[454] = 144'hfdc100c1fe8dfdd1fe9dff59ff1dfff900a8;
mem[455] = 144'hfdcaff33008bfe89016c012d0119fe61fed0;
mem[456] = 144'h011a0008fddefdc900f4fe5800bdff6eff4f;
mem[457] = 144'h01150166014601bdfe8a0098feaafe94fe3d;
mem[458] = 144'h0119fec2ff1afdf9017dffb50146fff2001a;
mem[459] = 144'h01b9ff67fe9600c2fe7afe64000700bc009e;
mem[460] = 144'hfeb6013201bcfe9c0002fe76ff14ff0e0117;
mem[461] = 144'hff1f008f00f8014801cbff32ffde0115fead;
mem[462] = 144'h0134008b00c8ffb3006700a4ff78fe4dfec6;
mem[463] = 144'hfeb40144fe9efe2800b4008afe8dffa7ff59;
mem[464] = 144'hffaf0442006c01e9ffaffc4202a20230028c;
mem[465] = 144'h003202ad0026020effa7002a01b7036b02b3;
mem[466] = 144'h01a802010123001afe21faf70316037a00b8;
mem[467] = 144'h00eb0215ff9e0105ff2dfdef001b043f03d6;
mem[468] = 144'h004d02d9016d001c015afdcb000b02c70055;
mem[469] = 144'hfe7dfd0ffd0e013d00cefed3febdf9e1fbae;
mem[470] = 144'h00c1022e0000ff1f0081fd4200b501a40134;
mem[471] = 144'h030d02f6ffebfd98fe0ffeda00d2fea4fefa;
mem[472] = 144'hff44021301ea02d3fee0fdd6ff7504890294;
mem[473] = 144'hfdc70337fe7effcdffc2ffe3003d03860112;
mem[474] = 144'h019f00e8ff8801ffff14ff1000520466015b;
mem[475] = 144'h013a006400e5fce1f87200cf00e6ff62fa4e;
mem[476] = 144'h01a000b402e6018dff5fff90ff690030ff23;
mem[477] = 144'hfe63fee9001a0009ffd0ff70016600290189;
mem[478] = 144'hfe9900e601cb0313019eff76ffda02b402d3;
mem[479] = 144'h007103e9021102760073fda402740267014c;
mem[480] = 144'hfec3fe0001f601b9ff19fe92ff3700dbffb6;
mem[481] = 144'h002cfff802d901e60223fe28ffbd00c8fe86;
mem[482] = 144'h0064021c01ac0125ffa5f96e00a0012efcb0;
mem[483] = 144'hff7a008901a80189025301fd012800050279;
mem[484] = 144'hfeb6ffd4026a035f015ffef3001304340099;
mem[485] = 144'hffedfe59ff3205d2ffec016dff02fd630381;
mem[486] = 144'h006fff4601d5010b02330088021c0295034a;
mem[487] = 144'hfeb40220031dffc5febd007d01620343fcf1;
mem[488] = 144'hfe7b01b60180008a0250ffafff3d0210ffdf;
mem[489] = 144'h009e00a1017601eb01bb008301ea005aff13;
mem[490] = 144'hfe3d016bfffd020400b6019f01c001740021;
mem[491] = 144'hffa2015404400109043502f70127008efcd0;
mem[492] = 144'hffc701df00d4ffd2fe4fff24ff1e019800cd;
mem[493] = 144'h010800420136ff4f00210030ffec0132ffa1;
mem[494] = 144'hffe6007b02760288fe0300d8005d0119ffd1;
mem[495] = 144'h01be01cdffc7012101bd00010128002d00d0;
mem[496] = 144'hff95fdfbff35ff61ff9401b3ff8c0056ff01;
mem[497] = 144'hff490021fe6e00ccfe3cfeb400a0fed9feef;
mem[498] = 144'h00e8fe48ffdd0065ffc40064007600fefdf1;
mem[499] = 144'hfec4ff0600f9ff75ff7bffe700e4fe83ff19;
mem[500] = 144'hffc7014b008a00820061ff94ff11ff26fdc7;
mem[501] = 144'hfdbf0151ffad0075fdfc007a002eff7bff51;
mem[502] = 144'hff4e0115ff47fea80137ff55fdc3ff89fe3e;
mem[503] = 144'hfe2fff01ff01ffcfff8eff67fe3a00890161;
mem[504] = 144'h0054fe8200f5fefe00340023002f000afe95;
mem[505] = 144'h002bfe3bff2bfdcc000eff75feb9ffb40245;
mem[506] = 144'hffd4fe7d008dfedbfe03016eff99fec7ffea;
mem[507] = 144'hfdd9fe99ff6900a5fea4ffd1ff47fe4dfee0;
mem[508] = 144'hffdbfe67ff11ffc4ffde00610006ff6f006d;
mem[509] = 144'h0153ffc2fed8011d016f00aa00eb015eff9d;
mem[510] = 144'hfe3afffd015401060067fe05ff4800f9fe1e;
mem[511] = 144'h00d80007ff44fda0ffdf0084fe4dffe3fdd3;
mem[512] = 144'hff3902310390ff5cfbd3fc2e00a7043603a1;
mem[513] = 144'hff4e0089004f0014f97efdbf010b02af03d3;
mem[514] = 144'hfe5d00760109fe9cfb89f8ae040c02fa0328;
mem[515] = 144'h0030ffcc0117ff40fbc3fcc9029803c204b5;
mem[516] = 144'h011c002c0398ffa7fb5bfe1a0184024d0451;
mem[517] = 144'h004efdfb0017067ffdaffd7cffd3fbacfa5b;
mem[518] = 144'hff8c002402f3ff07fe43fec502e7060105fe;
mem[519] = 144'h01e302f7037501adfdb9fd90031203ddffcb;
mem[520] = 144'hfe87ffd80314fd30fc12fca1028603a50394;
mem[521] = 144'hfd2100b2000200ecfbc2fac4fff8019c0445;
mem[522] = 144'hfd96008001a1ffc0fc1bfc7601dd04530380;
mem[523] = 144'hfe8000ca017ef656ff7f025202310178fe07;
mem[524] = 144'hffccff0a00a1016f00db008f00a001dc020c;
mem[525] = 144'h00f9017fff4cffdfff29fef100eaff9aff31;
mem[526] = 144'hff3a00580365feb0fc360030012f023601b6;
mem[527] = 144'h0065ff93026b005afd9dfe02030a01e3027b;
mem[528] = 144'hff5801080111fed1fcaa012c001201cb03f0;
mem[529] = 144'hfe5500d1ff80009afe2602b8ff3403970298;
mem[530] = 144'hfe7f01940352022e017c09d90231046901ae;
mem[531] = 144'h00b4fe4f009e01ecfedafffffe3503c9045e;
mem[532] = 144'h0147ff9103c301ce00190076fdb50456015f;
mem[533] = 144'h00bc0232feb4fd6efe7801d801d2fdaa00f6;
mem[534] = 144'hfe8f015803c70249008302b6031b027800ad;
mem[535] = 144'h00d6030102a8032806f604b90454012b012d;
mem[536] = 144'h0189fed6025c017e00fb0334ff050184049a;
mem[537] = 144'hfe6a014e01c0009afe7401a2fcd701a903d3;
mem[538] = 144'h003ffefd0249ff99021803740070013402c0;
mem[539] = 144'hff9b0048ff2ef858fab6ff78047404e9fff4;
mem[540] = 144'hfe99ff2afd9bfedaff62fe6501a5010c0188;
mem[541] = 144'h0163fe71001d00fa0010fe58019501210063;
mem[542] = 144'h001dff12fd44036c016c0191fd01fe1d0182;
mem[543] = 144'hfea9ffc40379ff510164027cff49042401aa;
mem[544] = 144'h00fc009ffe33fdfb001dfed0fefa003f003c;
mem[545] = 144'hfef2ff62ffa6ffd7fff60140fe95fde6fd9a;
mem[546] = 144'hff6cfe42ff7dfdaa0117fe58fea70021ffbf;
mem[547] = 144'h014efe1000e2fe7fff86fed3ffb8ff3bff2f;
mem[548] = 144'hfff400d80022fde800cfff92fdeefdc5fd99;
mem[549] = 144'h01400063fef200d5fef3012cfe44004efdd2;
mem[550] = 144'hfe36fffe0059fe6c00ca0024fe0cfe640044;
mem[551] = 144'h0136ff8eff9d0050ff63ff9efec4fe26ff15;
mem[552] = 144'hfee8ff13fe70007e0039fdc4015b0040fe03;
mem[553] = 144'hfddcfe51fe550012fe0afe5a00d6fe70004d;
mem[554] = 144'h0089fe7cfd99fe4b0121fe5900b80061ff6b;
mem[555] = 144'h00a800830111ffcafdc8ffc5011affbc0002;
mem[556] = 144'hff06fffd0155fe48fe3eff1c00ce00350120;
mem[557] = 144'h0103ff9b0159fe9cfe31ff31fe5301ae0179;
mem[558] = 144'hfe56fd9eff1afd9effd3fe1d00c0fe7efdbf;
mem[559] = 144'h010f0013fe07ffdefdfffea3febbfe12fe36;
mem[560] = 144'h011f014504a7031cfce2f75f034a00e303dc;
mem[561] = 144'h02ddffd403190018fe0efc8801baff9d0319;
mem[562] = 144'h01de031d03d200dffef8fab301a5ff760083;
mem[563] = 144'h0177ff2b01a9ff83fec8fb6f012401ef01be;
mem[564] = 144'h006cffbf02ca028c00c6ff3e022f00580125;
mem[565] = 144'hff3efc28f9cdfede0042ffc1ff0cf4f3ef12;
mem[566] = 144'h002901c9016d0312fe78fdfe0254016c027f;
mem[567] = 144'h00c0002c0387035a018dffaa0162ff3400dc;
mem[568] = 144'h0256024802330312fe6dfb5e012600c503dc;
mem[569] = 144'h01dcff5b02a60023fe64f81f0127fe81fe88;
mem[570] = 144'h01d9003803d802910309fcc70236026d0251;
mem[571] = 144'hfe38ff52fd20f7aaf659ff42ff77fe56fcba;
mem[572] = 144'h0176003602b201b9fe8bfebc0042fdeb002c;
mem[573] = 144'hffcf00e200fd019501d60102fe2afecfff42;
mem[574] = 144'h01cc026002ddff6afd6ffcd80304037403cb;
mem[575] = 144'h013300c90356032cffa6fad70072ff8f03a5;
mem[576] = 144'h01cf015f029d0126fe9df83f05d904070360;
mem[577] = 144'h000d02d901db023dff31fb0d045c04a2036e;
mem[578] = 144'h04de027001600104fc44f92c05470012fd58;
mem[579] = 144'hff82027702f3011efdb0fce9029602bb0476;
mem[580] = 144'h01ab01960402002401d6fec202ac00680134;
mem[581] = 144'hfebffbc3fb1d012a016f0001fd04f2f3f098;
mem[582] = 144'hffb8027504ba0342006afdf200fd029000ec;
mem[583] = 144'h0100034f01ec039203dd0003ffd2fedbfe98;
mem[584] = 144'hff5a00ef01c600e5ffcafbc40314030404da;
mem[585] = 144'hffd6023c01640145fcd0fd4404ad03ce0231;
mem[586] = 144'h02cd035304ac031a0264fe75046a03da01bc;
mem[587] = 144'h002c0096fcc2f897f3e4024c0157fd92f7c2;
mem[588] = 144'h00140025028401d1ffef00a10293fd8ffe72;
mem[589] = 144'h01affe5aff0b00a300190186006f01ddfff9;
mem[590] = 144'hffac03880251fe24fb1ef881035c04ce053a;
mem[591] = 144'h020903f5030a0223002afcd804b202ef02a2;
mem[592] = 144'h0143fdd8ff51002a004c00b3ff32ffecffb3;
mem[593] = 144'hfeb9fe1ffffefdfc011bfe23ff5fff71ffb8;
mem[594] = 144'h003b00e301ec00adfe970155fec4fffdff31;
mem[595] = 144'h008b0059012a00f600caffd5ffd0fde5ff31;
mem[596] = 144'h0175000c011f00c4fdf6010bfe3c0142fe21;
mem[597] = 144'h0176013d0087fde1fffb0106010aff26fedc;
mem[598] = 144'hff7c0135008400400089ffa0fea1feaf0123;
mem[599] = 144'h0127fdbfff5cfe0dfe6c0034fea9fdedfe5a;
mem[600] = 144'hfebf00b1fe31fdd5013e014c005200afffc0;
mem[601] = 144'hffabfec7fef9fee2ff6701be008fffeffdee;
mem[602] = 144'h0098fe79014601ee010d0074fed5fee9ff93;
mem[603] = 144'hff8400aaff50002400d9ff1600e900d4fe83;
mem[604] = 144'hfe74fe8201d3ff25ff70000b0036ff3effee;
mem[605] = 144'hfee0ffa7fff40116ff0b007100a70056ffe8;
mem[606] = 144'h00f70139fdf3ffaeffc8ff8bfe23fed0008e;
mem[607] = 144'hfe7eff7800acff39fe94ff84ff7c00fafee8;
mem[608] = 144'hfe51000ffec1fe8cfd9dfecdfe7401660180;
mem[609] = 144'hfddeff7f0003fd91ffe8fdedfe2a01dd0214;
mem[610] = 144'h00d901e5fff4ffb701f2034affab00f9ff9e;
mem[611] = 144'hfdd7ff5b0181feb3ff5bfe9c015600730072;
mem[612] = 144'h01b6002e005fff5aff0dfd30ffacff5e0161;
mem[613] = 144'h030c02dd0052fe020202007d045d019f054c;
mem[614] = 144'h00f9006900a6008e00ecfe150107ff31fef0;
mem[615] = 144'h00f800ef03060064024c026100be00ed0019;
mem[616] = 144'hffd4fe39fefe00e200e5fd3afe560322013b;
mem[617] = 144'hfe150093ff2800c5ff4ffdb0ff9800f9028b;
mem[618] = 144'hfde8fdf801f3fefc0022feb3fe1701e10174;
mem[619] = 144'h005301c2ff9dfd3bffba019fff4d025dfec5;
mem[620] = 144'hfe2b0099fe620097fe9cfe89ff13ffd9feff;
mem[621] = 144'hfeb6fff000d7ff2b00f1fef20164ff6bfe7c;
mem[622] = 144'h0048f6effdf200eb04f901fbfd8afdf900b2;
mem[623] = 144'hfe0101250228fed0ffa9fc3cfdcb0049018b;
mem[624] = 144'h014aff29ffd5fe3eff18006900effe6d00a5;
mem[625] = 144'hfe6fffc4fe0ffee3005bff4500b8ff5afec7;
mem[626] = 144'h02060091014600e0fd5e004101b800e10130;
mem[627] = 144'h011eff4eff07feedff65fe44008cff83ff57;
mem[628] = 144'h0160002c012e002101760161fe7bff7bffae;
mem[629] = 144'h0068ff8101d200f1ffec013cfe050024ff80;
mem[630] = 144'hffacfff10180ff50fee10142002400b900ae;
mem[631] = 144'h0145fe6fff98fee2007b002c016ffe630217;
mem[632] = 144'hfe5cfde3fffbfdd9008e008fff8efeeeffb1;
mem[633] = 144'hff740188fee9fe220110ff82ffd0ffde0136;
mem[634] = 144'h01ed0010feb4fe60ff09ff5f01c5ffd80047;
mem[635] = 144'hfea000e40014ffc6fe83fee3ffddffa6fe43;
mem[636] = 144'h001800f6ff1100dd0168ff43ff82fe9a001a;
mem[637] = 144'h005b0074ffc4011cffedfe2afe9cff28ff80;
mem[638] = 144'h0030ff9100abfe41fe9000080162ffeaff4e;
mem[639] = 144'h002eff7a012e0052ff45ffc3013b012a0020;
mem[640] = 144'h0480029d05170356fe4bf9d403d7fd760335;
mem[641] = 144'h01ab057403e1021ffdc2faaf032c0085007e;
mem[642] = 144'h045c03550150fde2fbd9f8ff002bfa5ff98e;
mem[643] = 144'h0231026f03d801fcfdc2004904beffa9001e;
mem[644] = 144'h03610433055f01330080014901a0ff91005a;
mem[645] = 144'hfee0faa0ff2105fcff4602d5fd8df7e0efa6;
mem[646] = 144'h020f02680438009bffe400e40033fe52fff4;
mem[647] = 144'h002701c2014afd94ff0c011afc11fd7cfa10;
mem[648] = 144'h03ac04c405f100b3ff70fc3700f801e00240;
mem[649] = 144'h019a040805a104de000cfd85056400e801eb;
mem[650] = 144'h02b004ef039000adfe8afe8901d40148fffa;
mem[651] = 144'hfed50000ff6bf6fafcc10299fdf2fb02fc11;
mem[652] = 144'hfecdffb001db00c2ff34ff8600e6fe5cfdfc;
mem[653] = 144'h005cfe76fea5fe76ff8e016fff6601ae0152;
mem[654] = 144'h0090049707ae036afd05fb67060a051303c7;
mem[655] = 144'h02ac0269040e017d0195fbe803cdfe99ffce;
mem[656] = 144'h01b20173006ffe67feb5ffa0ff23fdbf000e;
mem[657] = 144'hfeaa01950075004e0164feee0012febe0179;
mem[658] = 144'h01580009fde4fdd0ffe1ff87fed6ff99fdfc;
mem[659] = 144'hfe4201030169ffcaffb0fe44ff790027fed0;
mem[660] = 144'hfe61003afe9cff110154fe49ff6aff7afed8;
mem[661] = 144'h0160ff1bfe1cfe4200bf004efeeaffd80111;
mem[662] = 144'hfe9a002c00c7fe53fef3fe2a00cefdcbfe61;
mem[663] = 144'hfefbfec00055ff8fffc9fec4ff1ffeceff9b;
mem[664] = 144'hffec004f008effaffe9effc8ff80ff7eff5b;
mem[665] = 144'h0198ff0ffedcfdbe005a01e3fe9501d4ff45;
mem[666] = 144'h0019ff22fef9fdeefe96fe89fe7dfdb60155;
mem[667] = 144'h0113fdc0ff65019501c90096ff55005500bf;
mem[668] = 144'hfe29ff9e015e0047ff9a01a701be0146003c;
mem[669] = 144'h01090000fefd0087018dfedf008e01650176;
mem[670] = 144'hfec2ff0affdbff6aff95fdec010bff2200a9;
mem[671] = 144'h0126ff6b00a2ff4dfdb700aa011a00fa001f;
mem[672] = 144'h058600d7004effa1fd3afa38014c02fd038e;
mem[673] = 144'h01d70006fe6dfe32001dfba90487024b0168;
mem[674] = 144'h0579ffd3fddaff380121fc3efe40fe31fe48;
mem[675] = 144'h026f0030fde7ff43fdeffca504b8027e018d;
mem[676] = 144'h01b701e4ff99ff15ff63fe75031d01e8ffd8;
mem[677] = 144'hff6a011cff7bfe5100ef01f0fd7ef84bf60b;
mem[678] = 144'h0163029d00e90140ff8bfea60253009703e0;
mem[679] = 144'h00de03ef046a020c03180021fe5cfc2fff99;
mem[680] = 144'h01d701c3001dff8fff41fcae043b0221040c;
mem[681] = 144'h04c000e8fdf1fd80fd98fc3d027004250297;
mem[682] = 144'h058503370215009000a7ffd6031401550383;
mem[683] = 144'h027afde5fdcbfd7bffda01f7ffcafde4fb20;
mem[684] = 144'hfff6018f02370184004201acff8000dbfcef;
mem[685] = 144'h0057005401ca010500cbfef4fe6600a5ff9a;
mem[686] = 144'h0055ff93fcadfe03fd7cfe40072905f103a6;
mem[687] = 144'h027f00e80073fe740085fc7401dc00d20085;
mem[688] = 144'h010b012002af0130fdeaff43feddfdfb0071;
mem[689] = 144'hfec8022500e500360180fee7ffe9ff350186;
mem[690] = 144'h00f5ffe1ff590020fce5f5b5018c01f60035;
mem[691] = 144'h0216ff4f0067ff670082008c0142ff6f031e;
mem[692] = 144'h029ffeb500bbff8b01f6fdd4000e011a0130;
mem[693] = 144'hfff0012afd68029b00b10234004afc5df2d0;
mem[694] = 144'hff51fdb7002cfe79fcbcff4901d9026400f3;
mem[695] = 144'hfeaffce800dffe7dfda9fc1602340280024a;
mem[696] = 144'h0163ffba029600de0157fe11007e012601c6;
mem[697] = 144'hffecff5901a70022013ffe61ff3d0056fe3f;
mem[698] = 144'hff77fe4cfdff0262ff1efec1fef9ff28fe29;
mem[699] = 144'h00eb021a0258fe8cfd2c02c20044fe64fd52;
mem[700] = 144'hfec600f6ff4900ac015500d6fe96027eff2b;
mem[701] = 144'hfe5900b7ff66005e002201c000b3fe81ff61;
mem[702] = 144'h023c052a04a30276027d00a8037d00a102ec;
mem[703] = 144'hfeceff9d01ba019cff65fc9f0088002ffdcb;
mem[704] = 144'hfe9bfdfbfe34001e000501f2feeaffe9fecb;
mem[705] = 144'h00ecff61013001f2015ffdb90018feb6fe1d;
mem[706] = 144'hfe630064007f008ffd95ff8dfe9e02e5fd78;
mem[707] = 144'h01bbfe61ff90031cfecbff6bfe950297ffdc;
mem[708] = 144'hfda0fe63ff680321ff62ff30ffd300040079;
mem[709] = 144'h0067ff49fbe0008a02deff05fd56fb11fb6f;
mem[710] = 144'hfffefd5dfe260056ff0bfc26fff6003dfd69;
mem[711] = 144'hff50ff73ff35fed1fe59fdec004a01effd1f;
mem[712] = 144'h0002fe45fe0a0067003c002b000d0207ff2d;
mem[713] = 144'h00c1ff85fe32ffa800a1007dfe83fe81ff42;
mem[714] = 144'hfee8005d01780035fe4afd0cfffe0099fcfe;
mem[715] = 144'hfffdfe40fe41001dfb5b0089ff79008cff26;
mem[716] = 144'hff470029fe6a00e0febc00760227ffa700ef;
mem[717] = 144'h00ef00aa00bffee6fe60fe80011801b8ff3e;
mem[718] = 144'hfe2402550156015f013fff530058fe0bffda;
mem[719] = 144'hfe4effc200520109ff9ffed00099ff42006e;
mem[720] = 144'h0054ff3402cf00f2fda6fef3ff5f0011004e;
mem[721] = 144'hfee2fef9012100f2ff890196fe1c028402ad;
mem[722] = 144'hfeb901750328fecd043c094203c701b701e9;
mem[723] = 144'h0102fe06ffb800c6fe4e04b3fe140088012b;
mem[724] = 144'h005a0213019bff52ffb704f9fefa0142041c;
mem[725] = 144'h00e3010b01bcff91009b00f602d6024108de;
mem[726] = 144'h003901af012100520423046701ec02a802cd;
mem[727] = 144'h01f70102011e035f03f904b603c2011e019b;
mem[728] = 144'hfe65ff18ffa1ffafff58009a0162033103dd;
mem[729] = 144'hfe10fe4cff9e01b0011602930107008800f3;
mem[730] = 144'hfee2fecdfff001c0ff21023101840137017d;
mem[731] = 144'hff6b00b8027efaa402ea02800165056300b6;
mem[732] = 144'hff050024022cffbdffde00e4ff4a022d0200;
mem[733] = 144'h00be019c013bfef400effffe015900140089;
mem[734] = 144'hffbcfe97fe7a033ffe7e0064fc2fff03023d;
mem[735] = 144'h006b00690209013a00db01dfff26024a02d4;
mem[736] = 144'h014dff2fff09ff5ffe1f004c00c7fe97fe13;
mem[737] = 144'h012cfdc7fe9afddaff9cfec9feaafe3bff12;
mem[738] = 144'hffc801190167fe060163fe80ff0d01190020;
mem[739] = 144'hff69fe4100b4011fffb7ff8efed3ff5d009d;
mem[740] = 144'h0123fe2afe6efe8affecfe5dfdf20151fe95;
mem[741] = 144'h017a014e0038ff85ff5401770148fe53feb0;
mem[742] = 144'hfe35fe4900a40155ff0eff50fe1affc2fdeb;
mem[743] = 144'hfed000d5007f00c600ceffb1ff12fee400f6;
mem[744] = 144'hfe77ffde00edfe3600a80000014cff060061;
mem[745] = 144'h017700d2ff3400250119feb600fefe300069;
mem[746] = 144'h00fc007dfefcfdd20173ff860134fe76009f;
mem[747] = 144'hff6c004bfff9015bff37fe870022006c00d4;
mem[748] = 144'h00d70192ff77ff8dfe9e013d016601ac0112;
mem[749] = 144'h01df01bfff4900b80112007400b0fefa00d3;
mem[750] = 144'h0001ff9dff8dffc5ff39fe6eff91ff75feee;
mem[751] = 144'hfdfffddcfe57fdf2006cfec6ff5afeb90062;
mem[752] = 144'h0169049903350214020d02290204ffff0327;
mem[753] = 144'h020803c804a300c4ff11004cff820299fffb;
mem[754] = 144'h0234058603dafd3bfd9b0630fdf0fdc5fa9d;
mem[755] = 144'h01d701fa03e002b00115022fff4a00650081;
mem[756] = 144'h00410157044e01a2021c0267012b00f300cb;
mem[757] = 144'hffe3fbc2ff0502da004501cb000efa93000e;
mem[758] = 144'h004501f60142ffcdffc403c6012c00e9fe86;
mem[759] = 144'h025103040017fc490035019b0067ffe4fa28;
mem[760] = 144'h030b00db01b50170014effe6004903570205;
mem[761] = 144'h014702b0027e032a010501fc01cd019a00fe;
mem[762] = 144'h03760231033b023b0166014200c7015cfedc;
mem[763] = 144'hff8a0404007ff9dc00ed01ca0241002ffad4;
mem[764] = 144'h01c700b1020700a0feafff4400a7ffafff43;
mem[765] = 144'hffc6009c00f6feef0006006c01d6ff5d0078;
mem[766] = 144'hfeee02d4045c05ceff07ff5a0482035b024f;
mem[767] = 144'h01dd03c9027702ca010b02c5fef2ffaf0241;
mem[768] = 144'h037001e301d7ff340184fd1b007801c401dc;
mem[769] = 144'hffdb045200e6fe5e01a2fe7700f403b30242;
mem[770] = 144'h040700d4fe1bfc9bfe6efae7fed100ebfd7b;
mem[771] = 144'h001a026f0174006afded010a01cf02de021c;
mem[772] = 144'h011c03ed00eafee3fe220095000e01260048;
mem[773] = 144'h00bdfdcb02f7011aff680125fdfefd50016b;
mem[774] = 144'h00150267ff620026009f0134fedb01e40464;
mem[775] = 144'h022503dbffc6005f006700a2011bff23ff6e;
mem[776] = 144'h023201a6002dfe6700f8fedf02270352009c;
mem[777] = 144'h0044025100ea016f0106fe7000a6023c0245;
mem[778] = 144'h01fc01820273fe6700c600a2033d012f00d4;
mem[779] = 144'h0257013efe7200e704a1ff99fedd0070fa43;
mem[780] = 144'h010b02790262ff2201c401a300bf007700b7;
mem[781] = 144'h00a9fe5501c1ffab00d80151fe5bff6200f6;
mem[782] = 144'h0038032d036900c6fdfdffb5034f030f03d7;
mem[783] = 144'h018b048300cbfe350044fee6015f039001ae;
mem[784] = 144'hfe330004005003d0023702cffd7700760101;
mem[785] = 144'h00860191015300fb020d01e9fe9e006200e3;
mem[786] = 144'hfe0bfe7affc0015cff9dffc9fdac01c001cc;
mem[787] = 144'hffe2fea6fea702c1021effdffe00fec8ffe6;
mem[788] = 144'hff5a0049fe6703b501d0ffc9ff1afeed0008;
mem[789] = 144'h0100ff45ffe100b0020e010902e000b0fd18;
mem[790] = 144'h004c000c0193016c0122ff8b018a00cffde4;
mem[791] = 144'hffb1ffb200700018ffcefecf01ec021f00bd;
mem[792] = 144'hff5e00f0007001a702c40317ffe0ff3100ef;
mem[793] = 144'h01d2ffdd001d00fb02de007a0050fe2bfcc2;
mem[794] = 144'hff50002b019a038f023dfe270080fe0dfe2d;
mem[795] = 144'hfef0ff56065103f0ffbefff6feee03c603a3;
mem[796] = 144'h01a900eaff10014c00faff80008000d900b1;
mem[797] = 144'hfe4700bafea1fe390000014a01120013ff65;
mem[798] = 144'hff7903b5047102d8041b03f6fedffd95003b;
mem[799] = 144'hfe6bfe1201a1012a00ee012e001e00adfdf4;
mem[800] = 144'h0104fe4ffe26fea3fe28008fff6efeb6000c;
mem[801] = 144'hff6b013cfff3ff73ff7cfd5600a000b200e5;
mem[802] = 144'h00b601240087fdeaff7cffff008dff8cfdc6;
mem[803] = 144'hffdcfef6ff9afeab0025fe130118fe5dfe67;
mem[804] = 144'hfde20030fdffff24fe99007e0039fd43ff86;
mem[805] = 144'hff270109ff7dfdbbff980118008ffdbe001c;
mem[806] = 144'h00ccffdffee80008ff61fd62ff8efdd00051;
mem[807] = 144'hfd8bff78ffecfdb5fec4fe64fea9fda2fecc;
mem[808] = 144'h0153ffc300fb00bcfdfbfffb009bfe0dffc7;
mem[809] = 144'hff48001b00ecff2efd25012bffb8002a0078;
mem[810] = 144'h000bfdccff42013cfdbf0013ffc9fe71006a;
mem[811] = 144'hfd8fff8bfecb0150fdef013cfe5900f7fe46;
mem[812] = 144'hfe28fe2b014aff39015b0126008afe38fe91;
mem[813] = 144'hfec400fd00a20153009501a0ff38fee5011a;
mem[814] = 144'h0128fde9fda10096002dff9a0000feaefef0;
mem[815] = 144'hffa800cdffcbfe6efeadfde6ffccfe77ff2c;
mem[816] = 144'h055b037600affeacffcafd6e065a0082030e;
mem[817] = 144'h056200b20034fed800bbff5f046a011b019f;
mem[818] = 144'h04a500510081fe7afdc5f7a0030aff0affef;
mem[819] = 144'h0505028aff08fd4cfcdcfd35035f019501c2;
mem[820] = 144'h01cf036902290021fcd4ffc203e101220045;
mem[821] = 144'h007f0007063b02eaff5502b10077002cf97c;
mem[822] = 144'h010401cc009bfb16fec6fd890424ff300433;
mem[823] = 144'h03a400d70125fe2efe36ff86001afe7403a4;
mem[824] = 144'h032d015f0168fd200023ff8a04a302d6ffa8;
mem[825] = 144'h0208032ffe56fe0bff2dfcd405bb01b401e0;
mem[826] = 144'h04cc041b00ccff89feaefc1706500269015f;
mem[827] = 144'h027600fc0002fefb04de031300e1fbfb00aa;
mem[828] = 144'hffdb0094febdff6200ce01db0188008afe24;
mem[829] = 144'hfffcfe6201a1fe9afe24ffb1fee80087fe80;
mem[830] = 144'h01ee06cd015e01cf0117004e067706190176;
mem[831] = 144'h03b7027d0131fee6fcc8fdd002e50010015a;
mem[832] = 144'hfd43ff14ffe9fd85ff66020b020000a100fd;
mem[833] = 144'hfd2bfd11fcb1fd86feae02a8fdfd01ce018b;
mem[834] = 144'hfd64fc1401b1021902bffea4012b036006e3;
mem[835] = 144'hffe8fd94fecbff94ff1c02510015ff2a00c3;
mem[836] = 144'hfdefff72fdb5fef100e4024bff1701500048;
mem[837] = 144'h0023052b03a10306001a026d02ad07cc0886;
mem[838] = 144'hff1efd2aff650170011201db006b02de029b;
mem[839] = 144'hffaafebd00930395020700a30426020b04c1;
mem[840] = 144'h0093fe3c000e011201f9036cff88ff76000c;
mem[841] = 144'hfdfdfce4febb00db00da0358ff89fe84003c;
mem[842] = 144'hfd14fdb3fc3ffdcdfe7c02ecfee4031701c9;
mem[843] = 144'hff81ff59032e053801f7011e024302e4072e;
mem[844] = 144'h01cfffeafce5fe82fec600f7ff490028ff37;
mem[845] = 144'hfefffea3fe91ff4c01de00b3ffa4002201b2;
mem[846] = 144'h0192fd7efbd2ff8601df028bfc52fa2efd6e;
mem[847] = 144'hff00fd43fcf10136fea8029ffe0dffe2021a;
mem[848] = 144'h01520104fbd9fea4018f0480015403bf02e5;
mem[849] = 144'hfee802d0fd31fd670256033a003703bf0026;
mem[850] = 144'h0152026dfc8efe6f0107053002c300c702bb;
mem[851] = 144'hfe3801dcfde4fe50ff09ffef011400b900ae;
mem[852] = 144'hff1a0135ff53fe4bff5902bc023501960209;
mem[853] = 144'h01db05240555fb3a00bdfff5014908ef0d02;
mem[854] = 144'hff0601e9fce5fb2cff8cffa1004800d2044d;
mem[855] = 144'hfff1019efec6fe5b026502f402170070045c;
mem[856] = 144'h01260129fb7cfd97008504000017013100b6;
mem[857] = 144'h01d10203fcd3fcc1ffe0018400bf014a0166;
mem[858] = 144'h014f0171fd15fbdbff34033a012c02170188;
mem[859] = 144'h01c1fefdfe7b02520472ff810335025d0013;
mem[860] = 144'h009700fb00e6fe20ffb0fe6d00d9008d01f8;
mem[861] = 144'h005c00880067fea8011701b5fe8aff830173;
mem[862] = 144'hfdf500adfd4803430560043efcfcffed0033;
mem[863] = 144'h01220369fcd8fd79019d01b6003c022f023b;
mem[864] = 144'hfe48014d023a03ccff94fd27ff59fd740114;
mem[865] = 144'hffb5039d01f9014cff2900a0fe94fe7d0132;
mem[866] = 144'hfe5301af00a9009effbbff29fe4aff86027d;
mem[867] = 144'hffbc033e00ce02dfff37feccfe38004a0105;
mem[868] = 144'h0196013c01ac00bc01c4fe5100e4fe370172;
mem[869] = 144'hff6200ecffe50113002c0214016900a0feb2;
mem[870] = 144'hff96fff3011c01c801aafdd0ff92fded007c;
mem[871] = 144'h010d0293fecefddaff7aff4afdc3ff2902c9;
mem[872] = 144'h00bc0040038a02c10101fe040006ff23ffa0;
mem[873] = 144'hff27ffe603710374ffeafc70fccdfbfe0117;
mem[874] = 144'hfe6202bb0037009b02470200fd68fd58ff30;
mem[875] = 144'h01310018ff41feedff2cff97ff1200d0026f;
mem[876] = 144'h016aff8cff45003800670126fecc01b90312;
mem[877] = 144'h00cc00a7ffd40150feff0174018f0066fe43;
mem[878] = 144'hffd1003202b2ff5f0042febe00b9ffeb0243;
mem[879] = 144'h0058010a02ff01020132fe75fdfdff0cffee;
mem[880] = 144'h017304680360024401940063fcd4fdcbff09;
mem[881] = 144'hff1c046501a702bf0167feacfcd6fd60fe58;
mem[882] = 144'h01ed01bc0206fefefdcdfc44fd3efccffaf8;
mem[883] = 144'h01730358029003070328fe45008a007ffeec;
mem[884] = 144'h00bdff8703d50411023801c5fd62fe97feb8;
mem[885] = 144'h0048fd63fa5000d202fcffdbfe6efa33f378;
mem[886] = 144'hff4d02c8000203930059ff83ff50fe12fd86;
mem[887] = 144'h01b9fe39fea0ffb3fdfcffdffe75001afb24;
mem[888] = 144'hfec501ce039703c1019efd71fd23fe0fff09;
mem[889] = 144'hff4102e00282026003d0fed8ff52fcbaffd9;
mem[890] = 144'hff69024a01b804a604380274feb0fea6fc41;
mem[891] = 144'h006fff79fe67fea3faa0fd4afefbfd7afc19;
mem[892] = 144'h0164005c00e2010ffe9c019cfe49feb9018e;
mem[893] = 144'hff1e009b011b00490160fe3001c20147fe25;
mem[894] = 144'hff75056c02d6031600e4fcf9005e017a02cd;
mem[895] = 144'h019a027d017a03b801ecff31ff31001dfe11;
mem[896] = 144'hfd69fb77fd5cfe61fd8e018cfd58fe32ff2d;
mem[897] = 144'hfe51fc64fb82fdedfd7e0137fdb7fc9600d0;
mem[898] = 144'hfc93f932ff700006015405ddfc7200da08fa;
mem[899] = 144'hfe9bfcbcfd9efd5c00a200aa005cfc950385;
mem[900] = 144'h0174fef9fb60fcd2fef50003ffb2ffd101e2;
mem[901] = 144'h022c07cfff2afaa1fda5ff9b05ae04cef904;
mem[902] = 144'hfdf7fb34fbd700d102cf0442ff86ff35067c;
mem[903] = 144'hffa9ff02022b044a05d5060901ff036007c6;
mem[904] = 144'h0077fcc6fbf8ff6b00b2018bff5bfcb70332;
mem[905] = 144'h0014fb8cfafbfd6bfdffff88ffdbfd3002c5;
mem[906] = 144'hfdf9fc2cfa7afddffdb30092fea8fefc02a6;
mem[907] = 144'h00c2fc9101afff53ffe5001cfe3effc304e9;
mem[908] = 144'h01a100eaffacfe3b00dd003f01670180ff7e;
mem[909] = 144'h01bcfef4fede013cfe500053ff2101c80165;
mem[910] = 144'h02f5fefdfd53fe9002240068fd8ffd79fdd2;
mem[911] = 144'hffcdfa8bfd81ff6dfda9ffe1ffc9ffa70324;
mem[912] = 144'hfee5fdafffa20105fddafff9ff24ff99fe4d;
mem[913] = 144'hfeabfee00117fdd4008efe60ff84ff9bfdf0;
mem[914] = 144'hfe0bfdc400780022fe0dfda3011e00e9fead;
mem[915] = 144'hfda500fe00db004e00f7fe1bfed4fe81fe73;
mem[916] = 144'hff37fdde00f4fe150034ff86fe59fe69001e;
mem[917] = 144'hffbe00ddfe2afe94ff10fda3ffe3fdeafeaf;
mem[918] = 144'hff93fd7d0002006700ad010bfdc9ffed0069;
mem[919] = 144'hfda8fe8dfdc2fd8001040027fdc8fe45fda2;
mem[920] = 144'h00d1ff24003ffe6eff3fff9dfea4ffe800f9;
mem[921] = 144'h0110fd6f001bfe17ff8a0042fd9c008b00e5;
mem[922] = 144'hff57fe0dff82fd9c00610044fe0001220061;
mem[923] = 144'hfebc012e0125ff0c00bdfec00078012d004a;
mem[924] = 144'h0162009afeb8fe9a00a0fffcff690086fe2f;
mem[925] = 144'hffb2001dfedc005afeefffb0011cfef901b6;
mem[926] = 144'hff8a0076fdcffebc0047ff90ff10fd77ff10;
mem[927] = 144'h0015fdd6ffe0fe44ff00feb8fe5efe12fe5d;
mem[928] = 144'h002301aefe4bff32003c01cb01f30499013f;
mem[929] = 144'hfe57003400d8ff4702250236001e048001ca;
mem[930] = 144'hffa80208017cffbe023c02290343052dff73;
mem[931] = 144'h0004ff93ff590010ffd40234ff27028701b3;
mem[932] = 144'hfd82ff8900f5021b0070ff71feed02060317;
mem[933] = 144'h0062ff5ffd86fddc00570002ff16feff084c;
mem[934] = 144'h010b0042008d000e02ab003100ea05420002;
mem[935] = 144'h01bf01f6008f03e602e601f0008f03bdfcb9;
mem[936] = 144'h0059ff50fedb00f7ff9001d300800170011e;
mem[937] = 144'h000c006fff8b0212ff8601de002c028703a8;
mem[938] = 144'hfca70022014a00e9fecf02b5ff7a020e03dd;
mem[939] = 144'h01edff7bfed40194fba5fe8701250211fec4;
mem[940] = 144'hfebe01a8fe8d00820021019affe3000f0156;
mem[941] = 144'hffe801d50125fe8800c6012cff10ff1fffbc;
mem[942] = 144'hfeb6fe4ffd9201bdffea0018fc2afe73012f;
mem[943] = 144'hfdff001300690025008a024001360511020b;
mem[944] = 144'hff16fee4ffb0ff240109008500ecff0dfecd;
mem[945] = 144'hfe4400780043fe00fea800dcfdfdfe34000b;
mem[946] = 144'hfff5002000f30021fea0fec70088ff74fe88;
mem[947] = 144'hfeddfd9600b5fe47fe31fe3cfeaffff0ff5b;
mem[948] = 144'h00f3fdff00e4012700d5fdd9fe82fe4afee5;
mem[949] = 144'hfedffda100bb00d20006fdf0ff11fda100cc;
mem[950] = 144'hff15fd80ffefff5afed8fd6f010600e500aa;
mem[951] = 144'hfff00026ffb1fe17ff10fe18ff35fe8aff97;
mem[952] = 144'hfefdfe8ffe67fe330028003bfe10001efe7e;
mem[953] = 144'h006e00e8ffc1fff8fe69fda5ff2300e1fe91;
mem[954] = 144'hfdae001dfe3dfee2fe5cfef6ff19fe9400d0;
mem[955] = 144'hff8e0048fdebffdd008afe56fecefdb3feb3;
mem[956] = 144'hfe9fff24ff6d01bcfedffe26fe4e0156017a;
mem[957] = 144'hfe63ff6d0034fec400930164ffc7ff5001b8;
mem[958] = 144'hfd7a0068fec4ffeffe6bfe8efdbcfe560115;
mem[959] = 144'hfdd8fed9ff6afdfbfe4efe94fd8ffdf3ff60;
mem[960] = 144'h01140135ffe1ff8c000aff2200ccfdd1002d;
mem[961] = 144'hfddbfe39fde6010cfea500d2fdfdfe59000a;
mem[962] = 144'hfebeff12fe8b015c0094fe40fe380037fe4f;
mem[963] = 144'h00d90009fe820163feda0140fe48fdf6ff61;
mem[964] = 144'hfdd400f6017f00bcfe34febdfe1e00fffebf;
mem[965] = 144'h00bafe6dfee8fe5eff97ff9ffdd8ff2bffb9;
mem[966] = 144'hff94fde5fe13fe20ff62ff86016b0082008b;
mem[967] = 144'hff84ff400013ff45fed9fe490061ff19014f;
mem[968] = 144'h0135ffb7010b006300d4ff77fe6afe34ffe6;
mem[969] = 144'hfed5ffd0fee9fe4f015e01720030ffa0012f;
mem[970] = 144'h000cfe7fffab0067fe05fee6fdff0114fe67;
mem[971] = 144'hfebbfe50008401530017fe75005b000401be;
mem[972] = 144'hff81ff7200b4ff76fef300beff2bff5a008a;
mem[973] = 144'h00f7010ffecd01c40109febaff92ff660047;
mem[974] = 144'hff440161007aff51fe8dfeea000100b6fdc4;
mem[975] = 144'hfdfc0088fdd2004c006f013900b9ffaa00b7;
mem[976] = 144'hfed5fcad00110014fff9ffb0ff3ffcbefd0f;
mem[977] = 144'hfec3ff2a0082001cff930030029aff8ffdf5;
mem[978] = 144'h02bcfe9a0020fd6afedffe90ff9ffe33ff10;
mem[979] = 144'h00dffd450397fe5affd5fe87ff9afc98ff3b;
mem[980] = 144'h01aefea1028b00a3fe62fd3d001ffd6efcec;
mem[981] = 144'hfe83fe05fea20130009a0046fea2fe3701ba;
mem[982] = 144'hfec5ff39006dfff8fd40fdbbfd10ff760035;
mem[983] = 144'hff81fd38fff4fd9b007bfeabfe25fd20ffe6;
mem[984] = 144'hfe72feaa02cefd1cfeabfd4aff8efd7d001d;
mem[985] = 144'h000eff91027bffb4fffafef5ff18ffc5fe1d;
mem[986] = 144'h00acff8d0082ffb2ffe5fe3902bc0006fd0e;
mem[987] = 144'hff4efef300a5fd36018e007bfd09fe33008d;
mem[988] = 144'hffacff5aff45ff8e016500a1fe730098ffc8;
mem[989] = 144'hfe94018cfe4fff140015015eff91fed4fe8b;
mem[990] = 144'h00de018f01c8fde5fd55005000b6fce3ff61;
mem[991] = 144'hff34fd43fe4bfdb4fe99fcce02e50000fd63;
mem[992] = 144'h014401d9fedc02eb013301fcfe26fee1fe9c;
mem[993] = 144'h01c3015fffdb02ce01e7015d0116fcd6fceb;
mem[994] = 144'h0184000c00a1ffcefffefe4dfe74fe9dfd6c;
mem[995] = 144'h0446ffc1012a00f7fea60198021cfd5cfcba;
mem[996] = 144'h03efff7b0155fffeff9dfeaa013efdc1fcdb;
mem[997] = 144'h019d004200b905b10207004000270057010b;
mem[998] = 144'h0170fe0afe18fe84fdb1ffd8fde3fe1bfc53;
mem[999] = 144'h022dfe1eff4dfb3dfb6afc0affdaffc1fd1a;
mem[1000] = 144'h043800b1016cff3b032a01c200effd24ff2b;
mem[1001] = 144'h0316ffacffa30206005703d4ffe7ff9afedf;
mem[1002] = 144'h050bff3f000801360124fe030272fd5ffc04;
mem[1003] = 144'h0043ff32037106b4081300bdfdd4fe990208;
mem[1004] = 144'h01e1ffc202b9fe210072fe22ff3f000eff58;
mem[1005] = 144'hfe55fe36ff9cff4b001100e2011d01ac0138;
mem[1006] = 144'h01fa03fe02ffffa501040093056401430060;
mem[1007] = 144'h019dff56027bff7601cc02220149fddffcda;
mem[1008] = 144'h005500b10147fea1008a0084ff5d012e00de;
mem[1009] = 144'h00d9ff10013b019a004c0139fcdb00800272;
mem[1010] = 144'hfe18012802fe042103fa035fffc503760383;
mem[1011] = 144'hfe78fe7e0077ff3102ee01a8fda102f301ac;
mem[1012] = 144'h01a9ff7c0229ff6bffbe0009fd6702920269;
mem[1013] = 144'h03990351fc5df970002a03060334feb2fd74;
mem[1014] = 144'h011b008e031c034500a7035100a801d40098;
mem[1015] = 144'h0209014502f5059205a800eb00e4012a0163;
mem[1016] = 144'h012dffbbff19ffff000affee0062036903ac;
mem[1017] = 144'hfe7a0119ff7300f701a3ff96fb5201d3036d;
mem[1018] = 144'hff1c02400029ffa90259019cfd2b008a02b8;
mem[1019] = 144'h01ae0108fd5afc1afca6ff3e02d503d0fe35;
mem[1020] = 144'h004901b5ff38ffbf00b801cefec80070021d;
mem[1021] = 144'hfe53fe9901d8003efe3fff42ff6bfed5ff4b;
mem[1022] = 144'hfeddf9f0fc3d007a017e02b3fe0100dd04ae;
mem[1023] = 144'hfdbd009affc1ffcc0057fffffeaa027302e7;
end

always @ (posedge clk) begin
	q_a <= mem[addr_a];
end

always @ (posedge clk) begin
	q_b <= mem[addr_b];
end

endmodule