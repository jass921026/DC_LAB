`timescale 1ns/1ns

module wt_fc1_mem5 #(parameter ADDR_WIDTH = 11, DATA_WIDTH = 144, DEPTH = 1024) (
input wire clk,
input wire [ADDR_WIDTH-1:0] addr_a, 
input wire [ADDR_WIDTH-1:0] addr_b, 
output reg [DATA_WIDTH-1:0] q_a,
output reg [DATA_WIDTH-1:0] q_b
);

reg [DATA_WIDTH-1:0] mem [0:DEPTH-1];

initial begin
mem[0] = 144'h01e90026fb9aff71fc7cfd6e02b5041304be;
mem[1] = 144'h029f00c6fb58ffe4ff6e0094008c00effd3a;
mem[2] = 144'hf6ae0025fef4005c053107c8fd65fa86ff1b;
mem[3] = 144'h0505fbabf8bd01d9fbb3fbfa048a0881042a;
mem[4] = 144'h01a6019000fbfe7dfe40fadbfd32035a05cc;
mem[5] = 144'hfdf8fe9afe75fe25011f0013feb1ff42ffa0;
mem[6] = 144'h0208ff6efc140173fd32fdf002e40556019f;
mem[7] = 144'h038f0194fffd0169feabf99fff9802a3046b;
mem[8] = 144'h030c05a0fbcc0196fe6b00a0ff80ffd6ffaf;
mem[9] = 144'h034b03f5ff4900eefffafd95002203a502da;
mem[10] = 144'hf84afdb006adfc2d0437fd8afc4afe6e02c3;
mem[11] = 144'h011e00e8044cfdd800d0f573fc1f02ff064b;
mem[12] = 144'h00efffd4013e00b6ff53fcd004920a160392;
mem[13] = 144'hfd69f6bbf7e300c40191fdc8fbf1ff43fb35;
mem[14] = 144'h001afe7dfa16ff25ff1a0113035a03b8fcb3;
mem[15] = 144'h00c2021efec2003cfcc2fe01000502ff02f4;
mem[16] = 144'hff1dfeba00400103005dfefb012affd500c2;
mem[17] = 144'h001e005aff1cff2700bc00260014010401ae;
mem[18] = 144'hfffcfedfff14fe39ff59015f017600d60157;
mem[19] = 144'hffc6fe4eff5d0127fe06005b002b00dcfee7;
mem[20] = 144'h01e3010e006cfee6004bfdfdfe800175fe1f;
mem[21] = 144'h01cc01470051fe5601be0066ffb50151fedc;
mem[22] = 144'hfe15ffc2feaa003c014cff5d00a1fe56001c;
mem[23] = 144'h0021fdf70148006efeddfe0fff7b0122ffc7;
mem[24] = 144'h00b3ff50017efdfdfdc7ff53010e00480028;
mem[25] = 144'hfea4fe20017fff070002ff0afeaafe78ffae;
mem[26] = 144'hffe900d1fea70025001d00470145ff8800c4;
mem[27] = 144'hfefbfff0011dff6bffe4ff9900c9fea6ff7f;
mem[28] = 144'hff3b007500e5fe99ff26fe20008bff910060;
mem[29] = 144'h001a01bd00f601c801b7008afecdff7ffed4;
mem[30] = 144'hfe9ffe5afff0fe64ff8c0195ff4e01fa00dd;
mem[31] = 144'hff7cff02fe30ff84feb700f9feb9013a01ec;
mem[32] = 144'h00c001b4fe35ff4d01920115ff82fec0003e;
mem[33] = 144'h0191016cffb5003e00fdfe990003001900f8;
mem[34] = 144'hfecbff1c0031ff740150fea4ff0900a40183;
mem[35] = 144'hff4bffa800c8ff1201a2fe3afef2fe3a0023;
mem[36] = 144'hff9afdf30189ff2f005cfdddfeedfe57ff57;
mem[37] = 144'hfefaff98012ffe470196fe8afe4100a00159;
mem[38] = 144'hff61016701cafe36ff2ffe8e018e018501b3;
mem[39] = 144'h00f9feccff44fe21fed901c2feec017301cd;
mem[40] = 144'hfeb00014011bff20ffdb0045fe3200530190;
mem[41] = 144'hffbdfe94ffd9fe3300c1017efedaffe2fe70;
mem[42] = 144'hfeae00bb0067000400bf011600440165008e;
mem[43] = 144'hfe58fe8500c0010201a4016bffd200fbff17;
mem[44] = 144'hfe180097ff0a0183fe91015d007aff99001c;
mem[45] = 144'h00ee00c600deff8100ccff2cfe30010dffce;
mem[46] = 144'hfe52ffe9013dfed0009f00cf0042ffce00a1;
mem[47] = 144'hfe0ffffc0153ffc6fef2feca0073ffa8ffea;
mem[48] = 144'hff0b0091fe47fdba0117fe4dfefffd7f00bf;
mem[49] = 144'hfe3eff2efd7fff1e005afdbeff75008bfe18;
mem[50] = 144'hfddc00c7005a0025ffa900a6ff2ffdf4fe8a;
mem[51] = 144'hfeeefecaff17fec4ff130099fd87005a003f;
mem[52] = 144'hfec4ff7bff25ff18ff9afe010089010f0074;
mem[53] = 144'hfed3ff8a0124ff16011eff7dffbb005fff8d;
mem[54] = 144'hfe20fea0010dfdc9fdeffea700daff41fe11;
mem[55] = 144'hff82fef8fee9fde6fe69fd96008b002700ee;
mem[56] = 144'h00f60019fefcfe1dff12fe5efe2afd75fdea;
mem[57] = 144'hfd8dfec9ff17ffcdfd6600e3fda80057fd61;
mem[58] = 144'hfe510013ffadfea40095fec0fe4200c8fec0;
mem[59] = 144'h0063fdf0fdc1ff6cfdfd0041003fffb200ab;
mem[60] = 144'hfdda003cfe99fe3efe62fe96005bfd6ffecd;
mem[61] = 144'hff9bfdd4010eff72fdb5febfff02ff87fe46;
mem[62] = 144'hffc3009fff5dfebffdc4fe46fd58fde2ffec;
mem[63] = 144'hff9000d3ff20fdacff8dff48ff2dfe060011;
mem[64] = 144'h027204cf045800fe04e6018100d804460387;
mem[65] = 144'hffd0ff94ff5704bf0365ff82fdd0ff09fd25;
mem[66] = 144'hf581f993fff4011afbb4f907fba2f8beff79;
mem[67] = 144'h045406b701ba04310285fd3b011309480156;
mem[68] = 144'hfe82052904c8009f05c70594fcbfff0d033b;
mem[69] = 144'hff2cfffa002a01e8ff2bff0d0217002d01e1;
mem[70] = 144'hfd03037b0391031904d901cffe7503ba0205;
mem[71] = 144'hff8002dd0407fbfc0386044afde0000d004a;
mem[72] = 144'hfef202b6036e0438032e0157fe8dff8702ec;
mem[73] = 144'h0251047d04fe04ff031502a0fc8f018b01a4;
mem[74] = 144'hf999ff91fec8fd69fb3a02b6fcab00840253;
mem[75] = 144'h002f00c4016cff14ff4c0465fdde01ba045b;
mem[76] = 144'h03c10819033004150011f667037d0cf80213;
mem[77] = 144'hfe74f709fb03fcabf80cfd1efceafd9b01fe;
mem[78] = 144'h000500f7003f03b2025500a5fe3101cafd49;
mem[79] = 144'h00c8046b01bd019f04b7040efc37ffec0303;
mem[80] = 144'hff86001afe80ffbdfdc6ff8a00b200080074;
mem[81] = 144'hffe3fef7fe93ff99ff75ff2201410009fed2;
mem[82] = 144'hfeb4ff5fff8100ca00730102fefbff96ff5f;
mem[83] = 144'h01cfff690098fffa0063ffb8fe5afe78feb2;
mem[84] = 144'h0143fe3900adfeeffe3100c9ff04ff480093;
mem[85] = 144'hff3901a601a2ff42fe46ff6d00a60063ff4b;
mem[86] = 144'hfdef00130102013201420174ff8e01a0fefe;
mem[87] = 144'hfe3cffff007dff7c012e019e00f9fe860083;
mem[88] = 144'hfefdfe9a006f00d601b100990117016d009a;
mem[89] = 144'h001d0194ffdf000900f9ffe4fed700a2ff12;
mem[90] = 144'h006cffc2ff65ffec000c00a8fe8aff14fe5b;
mem[91] = 144'h008dff120087fffc01cdfeaffe0e00200210;
mem[92] = 144'h0084ffbd00a8ffc600ccfdc3fe8dfedfff68;
mem[93] = 144'hff2501470033ff84009c01410056febdfecd;
mem[94] = 144'hffc5002d0049008dff84fe48003aff69017b;
mem[95] = 144'h00eafecdfeb4fdee019f014afec9fed8ffa8;
mem[96] = 144'hfdc702b105df01a6007b0267f962fcca054b;
mem[97] = 144'hfb5201a9066400a3019a02b0fc780209020f;
mem[98] = 144'h0106049d0309029100e0fe5d0754ff0e0076;
mem[99] = 144'hfef8ff7b027d006101d30008f82aff720383;
mem[100] = 144'hfb90fde0035dfcdafeee0399fe78fba5ff83;
mem[101] = 144'h00caff9302e8028d0273010f014300680099;
mem[102] = 144'hfb52fd8f068901b602d002cffcd7feef03cd;
mem[103] = 144'hfe10ffe001c8fe04fe8f0090ffa2fb9a0011;
mem[104] = 144'hfccf02a908f700c7ffab0257fa9f000305c2;
mem[105] = 144'hfd40fcfe05a8009d00ea0358fca6fa3e03be;
mem[106] = 144'h021cffbbffe401fcfef00333062aff20fd56;
mem[107] = 144'hfe89fd8c0004022601230456038dfca1fea7;
mem[108] = 144'hfc10fdabfdf7038b0012ff5afc99fe46ffa6;
mem[109] = 144'h07fc0a160278fd18feb9fb150224ffed00bd;
mem[110] = 144'hfb2fff20065a001c023f0230fd1ffe59037d;
mem[111] = 144'hfe89fefb01ccff8302370272fa90faf902f7;
mem[112] = 144'hfe5ffea1017e0043ff58ffdf00b2011300ff;
mem[113] = 144'h0089019e015d006b015bfe2aff0afeb9fe92;
mem[114] = 144'hff2effa2008bff42feef00750042fe8afe16;
mem[115] = 144'hffcc0016ff520023fe3eff5d001afe950101;
mem[116] = 144'h0136015efe76fe6d01cbfe2e0065ff74015e;
mem[117] = 144'h0186ff26ff5901bc0079ff68009d000d0016;
mem[118] = 144'hfe75fe8bff480051fe7a00f5fdf702090095;
mem[119] = 144'hff90ff740009fff7004d0130010b0099fe24;
mem[120] = 144'hff4c01850093fdf5003bfdbc010cfe0eff52;
mem[121] = 144'hfff9fdeb00dcfe1a0150007bfe76feeb007f;
mem[122] = 144'hfe3b0073ffefffed0085fe8d01cf0031ff6d;
mem[123] = 144'h0089fe21002afe0c016b00dd0089ffed01e9;
mem[124] = 144'h01770000fea8feacfefcfe7e0081ff1000d9;
mem[125] = 144'h00a7fe4f00b9ffa1ffd0009701da00fbff3c;
mem[126] = 144'h01b501b100fc0103ffee01e9fec2005fff08;
mem[127] = 144'hfe49fed301e80146fe050162fe2dff540108;
mem[128] = 144'h000300560217052803d802a201e0023dfded;
mem[129] = 144'h041303e402ae031702d6fd4503dcff3f0359;
mem[130] = 144'h03dfffe800a900c0fe4bfc31fea40209009a;
mem[131] = 144'hfe5407e906c003e102130372033bfd5e0068;
mem[132] = 144'hfe58ff5d02d5034f03f904d501960356feea;
mem[133] = 144'h0026fd330063004e00a800e6008cfe31ff6c;
mem[134] = 144'h00ae022a0290038f037b00700067ff4502a4;
mem[135] = 144'hfcac01220280014502da021d00fa00bcffea;
mem[136] = 144'h014d0273ffa401bf0170009a0173ffba02d1;
mem[137] = 144'h014702d8007c0401023800a302c603450126;
mem[138] = 144'hfeaf03000000fe94fc7b012af6fe032700ca;
mem[139] = 144'hfbe6ff060246fe7c01540772fc40024eff57;
mem[140] = 144'h034f058f001000f1004f00ee0146fbc4fd19;
mem[141] = 144'hf8fa0030081a00c3fde802c9010004070207;
mem[142] = 144'h02bd041e038402f5001d003301e1fe6803c6;
mem[143] = 144'h0051037703f0033a01e002f30257022c01d6;
mem[144] = 144'h04200651020cfe03ff5bff9101a201a20129;
mem[145] = 144'h04cb0107fdc5fe0e0172013ffbe0fcc4f941;
mem[146] = 144'hfe7ffc43fec50042080b0781f9dfff5fff69;
mem[147] = 144'h0215ffa0fe8ffe6efbb2fef003aa033bfce5;
mem[148] = 144'h0689045f05da01cafec2fe79ffa0ffe500bf;
mem[149] = 144'h01a0030e000703b7034002ce037dff9efff3;
mem[150] = 144'h037b0368fe58fe5bfc91fec6fd3b01e0fa8b;
mem[151] = 144'h040c053102fd00e5ff1efe01ff18032affce;
mem[152] = 144'h04a7041d02a0fe51ffbcfd33fecafee5fe02;
mem[153] = 144'h050a048e03b3fe97fef5fd98fc49ff8efb77;
mem[154] = 144'hf8effbe8fef9fe71feb3ff61006902d600e3;
mem[155] = 144'h009603710202002bfcdcfae9fdf903b20266;
mem[156] = 144'hfe2bfbe801e0fd08ff50013d02de04010165;
mem[157] = 144'h02d1f871f977061b055b08140ba804ac0462;
mem[158] = 144'h039602b1ff66fe02ff45010bfd570024f8d2;
mem[159] = 144'h065705cd03cffe51ff06fc65fec5fdccfe34;
mem[160] = 144'hfe89002affcb020b02f40196fc92ff9dfb89;
mem[161] = 144'h013901cdfd9d01fd0383fc2a034502c80032;
mem[162] = 144'hfe780277006000f90063fee4069201c404aa;
mem[163] = 144'hfd02fca9008e025003f0fe2a0091fdb9f991;
mem[164] = 144'h02a00032fff000f003f204f7fc250258fcf5;
mem[165] = 144'hff88ff76ffe0febaff8bff9f03c1019a026c;
mem[166] = 144'hff6100cbfe7f00d7033dff6ffe50017ffce0;
mem[167] = 144'h016cffb9fd54fc80ff9502cefd70ffeffd64;
mem[168] = 144'h0068fe64ffa401b10549fc8403d1030aff6f;
mem[169] = 144'hfd770013ffd3039402bbffd8fd6805a0ff16;
mem[170] = 144'hfde001f9fee0018d0187087a0037ff6d0043;
mem[171] = 144'hfc9302cbff99004c0167088af8da0114005f;
mem[172] = 144'hfb8af71ffdc300a60574fa4c0729f899ffea;
mem[173] = 144'h05b505f205a3faf7f7d302b0ffc7fb9afe52;
mem[174] = 144'hfe36fefc017d011b035efe99fd3402a7fb82;
mem[175] = 144'hfefcfec5fe69028c030d01b6fbb70339febf;
mem[176] = 144'hff1b0097ff4a011effc4ffcc00a9022d01af;
mem[177] = 144'hffd20162fe8a0081ff9701b7009400ba0133;
mem[178] = 144'h017dffd30096ffba00f8020100d2ff36fe91;
mem[179] = 144'hfdee01d300870141fe350148ffbe0043fe1f;
mem[180] = 144'h0174fee6ff08022000f000760143fe380152;
mem[181] = 144'h00effe65ff1bff9200250120017301d3fe4f;
mem[182] = 144'hfe61fec7017a007a01ecff33fe89ff500044;
mem[183] = 144'h018000d5015b01e0008cfe71ffb6fe0dfede;
mem[184] = 144'hfe80ffe200bfffa00156ff44fe070133fe90;
mem[185] = 144'hff0bfde7013e00fb000e00acfdd4fffafe57;
mem[186] = 144'h009300f30025005afdca00aaffd2ffed014b;
mem[187] = 144'hff74ff7bff96ffa4ffb800fa0066fe1a0225;
mem[188] = 144'hfe120013ff6d003400d30077ffa60052fe02;
mem[189] = 144'hfe89fe3cfe94ff5aff6b00040021ff94feff;
mem[190] = 144'hfddbfe710166ffe600c5feab0160ff2effb2;
mem[191] = 144'hffc7fdcb01acff58016afe60010900c4feef;
mem[192] = 144'hff860117017d0188000d0087016601daffd0;
mem[193] = 144'hfdab0019fd5afe42017f00d5ffecfd2a0297;
mem[194] = 144'hff1cfb72fca3fd8a0073fe53005d002300bd;
mem[195] = 144'hffa5070e027d00e9023500b000c7059b01cf;
mem[196] = 144'hfef5ff04fffffeab00db03bd012301aa028f;
mem[197] = 144'hfe48fd51fdddfed4fe21008800b9fde10025;
mem[198] = 144'hfcd4010a00acff5a022e00bf0293fff404df;
mem[199] = 144'hfcb6007b0028fe8c004c01f1005effdc0311;
mem[200] = 144'h00d40205ff9dfd8001d6019002b800830393;
mem[201] = 144'hffcb020201e30092ffd002890287020fffa6;
mem[202] = 144'h01e700a4fe7efe21f901fe9bf7bf015501a0;
mem[203] = 144'hfdf3025b024fffdbfb970146fcd0007a00bc;
mem[204] = 144'h096c0d9c00ce0024ff75fc260127006cff6a;
mem[205] = 144'hf609fab5016c00d800abfdc0fa30ff4100b1;
mem[206] = 144'hffae03e900f30017ff30ff3f012eff8b04e4;
mem[207] = 144'hff6c009f0169feef0024000fffa302e00190;
mem[208] = 144'h01d8feaefdc7004401e4fe4b046d00b4fa90;
mem[209] = 144'h032e010dfa57037b001cfec600d6ff0bffdb;
mem[210] = 144'h014afe16ff4101ab02d8004dfc7f021801cd;
mem[211] = 144'h02530642039aff3d0138004a041804c1ffa1;
mem[212] = 144'h00c500c7ffc70390023cfe31004e03c30137;
mem[213] = 144'hff7200f90046fe57fe590183020a00830044;
mem[214] = 144'h03110055fd290004024c006401acff9bfc63;
mem[215] = 144'hff0c041101c2ffef0229ffdbff9b037f0034;
mem[216] = 144'h01b8fdc8fcb902d5ffb3ff0501ca0212ff60;
mem[217] = 144'h01b5024dff96035c02abffe1035100b3fe56;
mem[218] = 144'h057401a1014b02de02fa03250096034201f5;
mem[219] = 144'h04d1038500960353014e001dffac042a00c3;
mem[220] = 144'h06da07e306c8013a00b901e409780952022a;
mem[221] = 144'hf793fa820125ffa7fff8032bff6afc210087;
mem[222] = 144'h028b0190fdc6029effe3fcc00212002efadf;
mem[223] = 144'h032203b3010100ef01feff0002ca0361ff61;
mem[224] = 144'h07850363022f0096014fff230164028002b4;
mem[225] = 144'h001f012e0000fee1fef9fe0500000222f814;
mem[226] = 144'hfb58fcef0160fda2fe57010cfe7cfb64fea3;
mem[227] = 144'hffa6faaefc1f006dfeaffde500dc057afc78;
mem[228] = 144'h039404b70423fd700078fd02fe2f01ee02b2;
mem[229] = 144'h0114026aff8bff8a0096fea200a4feeb0028;
mem[230] = 144'h03bdff8a0268002bfcaafea7fee50284fb65;
mem[231] = 144'h039700a502f3ff26fe94fd6a00a0032301a7;
mem[232] = 144'hffca04e102eefa88fd5cfe4fff000154fd9a;
mem[233] = 144'h039d050e0400fefffeeefc01fd6cffabfc14;
mem[234] = 144'hf1f2fcdcfff5ffabfecaffbbfc0ffebb0275;
mem[235] = 144'hfc7c018f04d7ffc3fd0ffd72fc4301ed02c8;
mem[236] = 144'hf5abf6e7ff5b0013fd2afd24fe6701c6fdbe;
mem[237] = 144'h0df90023f9fa059806c004ef065005ac050e;
mem[238] = 144'h009301f00192fe18ff2dfd00005002eef8ac;
mem[239] = 144'h02d8026c0257ff1dfd0afb87ffdd020dfdda;
mem[240] = 144'hffac0114006701b003b404dcfb6cfd8002f6;
mem[241] = 144'hfddd02820617072d02610264fda102d40402;
mem[242] = 144'h003e0600041701d8fbbef82c047b03d0ff62;
mem[243] = 144'h00c4fd470045061403cc0661fadffba202b0;
mem[244] = 144'hfde300ba006bffb2047e070302dffb02011d;
mem[245] = 144'hffc8fff6ff1dff090034ff48016503860233;
mem[246] = 144'h01a8fde10140065c03e306fcfcc9fca60240;
mem[247] = 144'h01ac0112ff84fe8a0429061f0131fa4501cb;
mem[248] = 144'hfcf7fe2803bc0748035a0169fd00036602d8;
mem[249] = 144'hff52fd4c009b036102c50754fe28fcee04d4;
mem[250] = 144'h04c40155fffe02a4059c03130712fe36ff0b;
mem[251] = 144'h00aa015dff74048105d209e202e3fd6dffc8;
mem[252] = 144'h01eaf78afcfe076703d60486fae9fe200342;
mem[253] = 144'h02a609f005acf660f168f9b401d4fceafd6e;
mem[254] = 144'hfda5ff2d047e0420013a044efd0dfe530395;
mem[255] = 144'h00effd5d022505fd047b0652fd82fe110343;
mem[256] = 144'hfd5fffb100dbffc0ff42026efe89fcc2fe0f;
mem[257] = 144'h007a0064059affe00127069b00ad0126014b;
mem[258] = 144'h04c5067f03a6fe18004d031703db073dfe54;
mem[259] = 144'hfce3fca7025b023900af055efa69f47efce0;
mem[260] = 144'hfdadfe81fd84fe5affe501be043dfe94fb7e;
mem[261] = 144'hff67006dfeb101fd013b01b300300045ff93;
mem[262] = 144'h007d002401a10148fd8a0545feedfc02ff49;
mem[263] = 144'h018bfebaff3e0220ffcd004a056bff54ffd3;
mem[264] = 144'hfddbfe4402b0fbb2012806d302b7fe5fff75;
mem[265] = 144'hfebafc920007fd2bfe6703760407fee5fd4e;
mem[266] = 144'h012cffe3fdf6024affe8fb31ff8f0191fe35;
mem[267] = 144'hff39fdd9fe2a01b600e4fe0f01bafb4afcd6;
mem[268] = 144'hfb2af604fd0b0097011907a7f10ef171fb53;
mem[269] = 144'h03ff097f06f00077000efdce035104790335;
mem[270] = 144'h008dffe703e30084fdce05f401f4fec402cf;
mem[271] = 144'h008dfe87011effa0fee703fb03dbfe30fdde;
mem[272] = 144'hffc2fd79010e00db019dffedf942fcbe02ce;
mem[273] = 144'hfd030068072401cb0049fc8aff86045e0469;
mem[274] = 144'h00d308ea03ae0097fdeeff410a4601620027;
mem[275] = 144'hfb06f75c000201590302ff37f932f8fcfe5c;
mem[276] = 144'hfffdfd78fd6cfdeeff6b010aff40fc1c00f7;
mem[277] = 144'h0132030e011b00edff8cff1100b300bc0163;
mem[278] = 144'hfc8bfbca03d30023009b0169fa7801fe0229;
mem[279] = 144'h0280fe84fda4fdf500d0012bfdbffaaa011a;
mem[280] = 144'hfa88001d060200e7030ffc5cfe3c044f039b;
mem[281] = 144'hfb13fc6b02e5ff74034900e2fb5cffa602b3;
mem[282] = 144'hffd8004dff05ffc803ad03f60401fa12fe09;
mem[283] = 144'hfe86fcb9fc41026d04ab058300ddfbd6ff0e;
mem[284] = 144'hf8dcf280fc7203b400d9004c00b9fbc60154;
mem[285] = 144'h0c0e0bd70515fd68fb66fc860408feeafe9f;
mem[286] = 144'hfacbfe9403df02bcffe6ffecfb3701ce020f;
mem[287] = 144'hfdb0fddfff22ff5103110155fb10ffbe0260;
mem[288] = 144'h0221020e05faff670309029d03a6feba0078;
mem[289] = 144'hff6100da06dd00ddffea04b10540fec6fb94;
mem[290] = 144'hfc7f018e0257fe50fb4901ba02d30146fee4;
mem[291] = 144'hfeab052b05d4012e033105eefd6afdcafe27;
mem[292] = 144'hfe6000bb042bfd6e021506600602006dfcce;
mem[293] = 144'h002afdf5fe9c0155fe9801a2014a00df01e1;
mem[294] = 144'h001501ed03e4001e03450550037201f0fedb;
mem[295] = 144'h00be01e60093ff63017901b602c7ffc3fd98;
mem[296] = 144'hfedb0007046600c601b506f30609ffc9faf0;
mem[297] = 144'h0077038604dbff2103370719043bfe80fc0d;
mem[298] = 144'hff0fff0bfe6f0083ff43fb7ffdca02d9ffd0;
mem[299] = 144'hfe3102a3ff3e0216fff902b702b90396feee;
mem[300] = 144'hff440303fe2f013a032a0300f3b6fa44fc14;
mem[301] = 144'h037504410521fc49fbf0fbaefd2002b205cf;
mem[302] = 144'h005402a006a50246ff80053d0447ff39ff39;
mem[303] = 144'h01b3015a0471fff8018606eb02e30207fbf4;
mem[304] = 144'h011a000bfe5100bfff630054fee4fdd8fe19;
mem[305] = 144'h017bfe44001dfdb6fdff0145fe4500860030;
mem[306] = 144'hff6efe94014ffed70100fee6005100aeffaa;
mem[307] = 144'hfe24003b002f00300144feaefe540101fed7;
mem[308] = 144'hff8800f3fed8007afe7eff8fff3affe7ffe9;
mem[309] = 144'h0143007a015f0153000200e200dd01a50058;
mem[310] = 144'hfdddfe56fefb0083009efff90049febb00c9;
mem[311] = 144'hff32fe21ff9b0164fe97008bfe8a00850019;
mem[312] = 144'h006ffe100097fe04fef600de004a00a40030;
mem[313] = 144'hff3f0070012bfdd2fe9efe24fe85fe2e0033;
mem[314] = 144'hff0eff40ff7b00d5ff79001e012c0059006d;
mem[315] = 144'h0067fe1eff41fed3018c0054ff540073ff00;
mem[316] = 144'hfe5dfe40fed900bfff77ff43015c001a0166;
mem[317] = 144'h00c5ff53fede0136feb4fe6300cdfe9e002a;
mem[318] = 144'h0096ff9c009bfe19fef2007b0000fde0ff50;
mem[319] = 144'hffc2ff19fe060107ffe0fecffebffecbfdd0;
mem[320] = 144'h00cbfe03fd66ff0201b4016503b3019ffecc;
mem[321] = 144'h0242fe84fb4402ec032b006bff670094ffd5;
mem[322] = 144'hff0eff59fe1403bd0434fe39fcceff3802a7;
mem[323] = 144'h05de04c2ffc8ff07023e03a8065403ac0453;
mem[324] = 144'h00a000edfdbc0113ff480356024a023a02de;
mem[325] = 144'h0069ffadff390009008600be013dff68ffea;
mem[326] = 144'h040d0258fd68006d03cd046e02d9ff7c01b8;
mem[327] = 144'h00e0ffc0ff05ff6e02280285ffb6ffd10113;
mem[328] = 144'h0338ffc6fb90059b062803ab021800a603a1;
mem[329] = 144'h023c032dff1f03f40334047effd501bf01cb;
mem[330] = 144'h0907062f00ffff4c02ff03b605e601fe013c;
mem[331] = 144'h070303a9017d00cc02fb0319037e02290228;
mem[332] = 144'h0b9206a50516011704c9017f056605a605ea;
mem[333] = 144'hf52af828fe03f770f47bf9eafed0fa97f739;
mem[334] = 144'h0106012afd1404b402ba018000e100f700c9;
mem[335] = 144'h027600dcfe4e038b02ac047b00e3030500ce;
mem[336] = 144'hfcd500ae02b602d001e5049e0302fea5fca6;
mem[337] = 144'hfdb2ff7600c7031101530120009e005c0394;
mem[338] = 144'h03a1ff59fdd300defcb0f9e203b205730461;
mem[339] = 144'h011c074308d200a002a30273006efea7fd3d;
mem[340] = 144'hfabafed500280119042f036000b4016efe43;
mem[341] = 144'h016700bcfe5c000cff5bfe8affd8004800d1;
mem[342] = 144'hfddd02c502060061042802d201ae007b0376;
mem[343] = 144'hfc130010010a00d4039c0385024900d4fe1c;
mem[344] = 144'hff0cfce800c800ff032e03d3019c00630210;
mem[345] = 144'hfe85fe8b011d014802b904fd02ba006aff59;
mem[346] = 144'h05ed024efd74ff05fd810229fb67048000b1;
mem[347] = 144'h0027ff8000a602a9ff2e0743fec2ff59ff20;
mem[348] = 144'h0659092902b100fc0413ffadff26f855fb63;
mem[349] = 144'hf9a205da09d2fc8ffc9c012dfb65fefd01cb;
mem[350] = 144'hfe1b02e60358034602e802e00166fe64052b;
mem[351] = 144'hfcee00d0000002e2011f01ec01a201a8ff1a;
mem[352] = 144'h00c30368008afc77fe68fcdcfffc015efdd2;
mem[353] = 144'h023aff30fd2afff500ffffb7febefa72fee7;
mem[354] = 144'h024ffc77fe9f0319091807befcaaff89031c;
mem[355] = 144'h05c503230035fa76fdebfe8b012cfe92ff97;
mem[356] = 144'hfeeb010bff61feebfda5ff61fbe0fee5fde6;
mem[357] = 144'h0283ff7c01abfd6bfffa02bdff8f0111ffe0;
mem[358] = 144'h01670288fc8cfd7cfefdffa7fffafd3dfb22;
mem[359] = 144'hff0c00670020ff40fc2301fcfeaaff51fc44;
mem[360] = 144'h02d401ddff6cff6e031f0086fcb4fcbe001f;
mem[361] = 144'hff7902a7fff6fc020022006cfeabfda5ff1f;
mem[362] = 144'h008002840000ffddfc4b0071038905380140;
mem[363] = 144'hfd9101bdfffe01c6fc1bffef005f019ffe84;
mem[364] = 144'h09a3099a027f002f03c2fc84036907e2056d;
mem[365] = 144'hfc6ffe50ffae014b003d02ca03450159fe96;
mem[366] = 144'h019303edfe5bfad5ffcc0041ff91fb5dfde3;
mem[367] = 144'h001600330182fc100106ffde0069fe79fd90;
mem[368] = 144'h0058fe570098fee4ff31010a015ffe630127;
mem[369] = 144'hff4c0057ff0efe9dfeaaffcd011401750179;
mem[370] = 144'hfe49ffd5fde7fe53ffc30140fdf900ee0029;
mem[371] = 144'hff5700b00078ff2700dc01d200aa0074fff7;
mem[372] = 144'h015601c00171fe7600ce00a0ff470101ff08;
mem[373] = 144'h01310002ffc300dc00660112007a008dfe72;
mem[374] = 144'hff820165ffbafefe000b00a6007bffe200a2;
mem[375] = 144'h00b1feadfef6ff6cff63ff8a012800ec0047;
mem[376] = 144'h015cffc0fe49ff14fe40016e00a0fed8ff00;
mem[377] = 144'h018d009c000101760174ff54fe5cffc500a4;
mem[378] = 144'h00df00a2017d0007fe48ff81008500da01db;
mem[379] = 144'hfdc8fed3fea9ffb3fe5a00bc0064fe9800c3;
mem[380] = 144'hffb6006cfebffdf3fecafe66ff49ffdb0115;
mem[381] = 144'h01c8fff9ff1501d3ffc90114018d00770081;
mem[382] = 144'hfec7fff9fedfff1ffe2400bd0002ffcb006f;
mem[383] = 144'h001bfe7ffeb00081ff13013e011dffafffc2;
mem[384] = 144'hff470096009601dcff6d0024ff1cfdbefed2;
mem[385] = 144'hff00fe77002e0162013efcf4ffcbff86007d;
mem[386] = 144'hfeecff1fff890010fe43003b005bfe80ff07;
mem[387] = 144'hfdf9fdb9fdf1feb0fdfefe23ff64fe4bfe94;
mem[388] = 144'hff0aff5dfe5d024cfffa00fd0051fdafffd4;
mem[389] = 144'h00fcfe5100ba00c300a5016700ceff8cfe67;
mem[390] = 144'hff52003dfd4d009afeadff47fe800084fe16;
mem[391] = 144'h0033fe39fe87ffb600ae00450067ffebff22;
mem[392] = 144'hfd9cfec0fe8302abfef3006efea0fd6afffa;
mem[393] = 144'h0002001cfdf202b4002d002ffe82ff8affe5;
mem[394] = 144'hfe0c005cff0fffdeff6c00a7fda0fe94002a;
mem[395] = 144'h000e006dfdf9fe04015700b1fd8700cc0009;
mem[396] = 144'hff43fdcafe960002fd46fe5c00a5008cff9d;
mem[397] = 144'hff66ff2dfe2efcee008fff5b01180099ff62;
mem[398] = 144'h0077fda2fec501590032fe55fe5a006dfd62;
mem[399] = 144'hfdf800e300e700ccfe20ffec006d00a3ff26;
mem[400] = 144'hfe7a00710010fcbdfd26fcea02cd01d4fc0b;
mem[401] = 144'h051102bcff7efec3025bfecc02a1fd08fe70;
mem[402] = 144'h048100f100510556091602fdfed0fff802b6;
mem[403] = 144'hffd804300260fc87011effb103dd020cff32;
mem[404] = 144'hff6c000100eb00aefdcdfe57fd5b01fefe33;
mem[405] = 144'hfef700b4fefa00d1fe9a0124015c035b016f;
mem[406] = 144'h0026025dfed9fe4e0139fde9016400bcfbdb;
mem[407] = 144'hff250053022e00000031ff39005d02edfc61;
mem[408] = 144'h01cffeedff34011d0053010aff28fd62fe17;
mem[409] = 144'h032f033101eaff3700bbfd9ffdd500ecfc66;
mem[410] = 144'h009f02edfe73008f006105cc032302c400eb;
mem[411] = 144'h006901bd01abfff8fc08fee1007003b4ffcd;
mem[412] = 144'h07a0058f046501160133fef704d303410272;
mem[413] = 144'hfa4afaf3ff07ff21fffa050e00efff080412;
mem[414] = 144'h02c703880010fd9500c4fe08021d0011fc8c;
mem[415] = 144'h021900430027fd5a00f7fd9b01db0204faf3;
mem[416] = 144'hfdcffcc9ffd2fe31fdaefcc4ff44ff39fecc;
mem[417] = 144'hfca300c7ff1afd7ffca8ff0c0240ffa40092;
mem[418] = 144'hff8efeeafd53fc31fe20016e00940042ff91;
mem[419] = 144'hfbdffe3200c400d3feb3fd9afd5afe4dfdfd;
mem[420] = 144'hff13fe4cfd77fde0fd44fc77ff3afe45fe71;
mem[421] = 144'hfebfff4c000e01a9ff9a002500a9fed1fe98;
mem[422] = 144'hfec9ff3fff39ff70fdbafcf80166fe9ffef3;
mem[423] = 144'hfdf0fff60074fcf6fd26fbc7fe980107fe51;
mem[424] = 144'hfd24fea200b3fc2afe10fdcf01afff4ffe5a;
mem[425] = 144'hfb5dfe74009cfd10fe8cfccbfe25fd6ffe00;
mem[426] = 144'hfda9fcf3ffb8fe15fe7ffd25fe78fe5bfd89;
mem[427] = 144'hfbe4fd62ff97fd400137fe45fcf4fe17ff47;
mem[428] = 144'hfd67fd2afca2fd6fff03011dfc69fd78fdd2;
mem[429] = 144'h022dfdcfff04feb8fe09fc76fb9cfdc7ffb7;
mem[430] = 144'hfe3bfe4fff13fd18fd1afd96013efe33ffc2;
mem[431] = 144'hff03ff6cfdd9fef0fffafdcc00bffdb500ed;
mem[432] = 144'hfe5700c10012ffb10110fdd0007b007afef8;
mem[433] = 144'hfe87ff7601b600cf0011004e00fb0122002d;
mem[434] = 144'hfee000cdffc900c6ff6400c9fec600cd00a8;
mem[435] = 144'h009bfeac0023015fff9efea4ff0effc2012a;
mem[436] = 144'h00ab00de0098fec000d0ff790154fe36fe62;
mem[437] = 144'h0022012bff3f0196fe4400caff12ff05ff64;
mem[438] = 144'hff6b0100ffc8fddefeeb0244fecf01150138;
mem[439] = 144'h01a3ff41fe0fff33004400a600b6fdbf00da;
mem[440] = 144'hfe0d0165fe7bffc6008e016b00d3fe3effbf;
mem[441] = 144'hffacfe19ff77feac015001f8fe8a019cfede;
mem[442] = 144'h0026004dfe5d0007fe6fffdc00e8fee6fdcd;
mem[443] = 144'h01b6ffb6ff550095014700f10099009dfdc1;
mem[444] = 144'hfe0efe39fe1a012bff97fe9f00eb0062fe32;
mem[445] = 144'hfe81ff1eff07ffabfdaf0137017400a2fead;
mem[446] = 144'h0059ff110058fe2bfdf3ff14016b00befed5;
mem[447] = 144'h00faff59fe02feaefea5ff48fef701d2fdf9;
mem[448] = 144'h00b1ffea01510091ff13fdcdff5600b90104;
mem[449] = 144'h01f9fe3cfeb8ff0900d00189fe72ff9afee2;
mem[450] = 144'hfec4011b0146021fffb600ad00c201effe89;
mem[451] = 144'hffbd00c10092008c005500c5017300060063;
mem[452] = 144'hfe2d0058febbfe16feaa00daff22003d0167;
mem[453] = 144'hfe89fe3201100080ff5800e8004a0087fe36;
mem[454] = 144'h01cfffa60075007ffe1cff40ffc6fe82ff0b;
mem[455] = 144'hff36ffed00c70131003bfe7d017bfe92fe19;
mem[456] = 144'hfdd5ff4cfdd2fdd200e3fdf1016fff97fe9a;
mem[457] = 144'hfdbffdf9ff6a00a7ffe4ff06fe8c0090ff48;
mem[458] = 144'hff5c00c7fddc00b500f6fe9900e600d0feab;
mem[459] = 144'hfea20008010efe1800b2ff17003b0100fdd5;
mem[460] = 144'h00defdd300a400fbffde008f0010ffb1ff9b;
mem[461] = 144'hff03fde70032022a00c0014400c60020008b;
mem[462] = 144'h01c6ff9ffe67fe760040ff400017fe7ffedb;
mem[463] = 144'hfe7dff4bfdc8fe1efeaf000cfeb30000fe90;
mem[464] = 144'hff4700cefc58fd2fff2cfcdbffbb042b00c0;
mem[465] = 144'hfbecfe85fc58f9c7fbe9faed031802840127;
mem[466] = 144'hfb69fe3ffed6fbfafdfe010f02d9fe2200ea;
mem[467] = 144'hfcddfcc0fbacfcc9fdd3f90c02e70574004f;
mem[468] = 144'h0059ffadff92006efc94fda4fd85002a04fd;
mem[469] = 144'h00db017500790197ff7f0062ffbbfe70fd65;
mem[470] = 144'hff0dfff6fe1bfbbffd80fd5f010502edfef9;
mem[471] = 144'h00aefee9010d005efce6fcb8fc73ff710255;
mem[472] = 144'h004a024bfb2ff9dffcaffce20330028103d3;
mem[473] = 144'h00e8fec8fff5fa28fd5bfbf6ff5501d800e1;
mem[474] = 144'hfafdffa70023fe23fef90223fb4afb840151;
mem[475] = 144'hfeebfc8d0089fce1fdfcff01fb7000e603e6;
mem[476] = 144'hfa9101330150fccdfefcfe5707b30379001f;
mem[477] = 144'h031cfb06fd2607820839032cf99bfee0feea;
mem[478] = 144'hfd38ffadfec7fbbffc7efbee022302c300dc;
mem[479] = 144'hfdeb00acfd95fba0fc7cf9d3fe6902910106;
mem[480] = 144'h001a01d4fa24fe2cfdfdfeb803c8fec1fef8;
mem[481] = 144'hffb2fb51f75cfcf7f941ffb6ffd6fb5303c7;
mem[482] = 144'hfe4efae6fd51febbfe820265fbc5005102f5;
mem[483] = 144'h016cff6ffe7effc9fd39fe9b053304170109;
mem[484] = 144'h02c600deffc20021fec8fd68fea7ffb4009e;
mem[485] = 144'hfea70015009f0135ffafffa8fdb8ff96ff19;
mem[486] = 144'h0134fec1f99efdcbfc84fb940419fd1bfdec;
mem[487] = 144'hfea1027b0153008cff62f9d2018c003cfebb;
mem[488] = 144'h024bfe3afa01fa5dfc76ffb7ff34fc39033f;
mem[489] = 144'hfff9ff64fda5fc1bfaeafb3fffd1fdc7fd1a;
mem[490] = 144'h02e0033e01b00202fe2cfd360026026f00a5;
mem[491] = 144'h009a02d8012b01b9fd6df8bb030e0480016a;
mem[492] = 144'h040d06910222fdc3fd7dfeab04a4091802c3;
mem[493] = 144'hfc2dfaa2fd1706c908aeff69fc2afe15fc12;
mem[494] = 144'h0073fddaf9fcfd91fcadfc5b012dfc76fed7;
mem[495] = 144'h009001fdfaf3ff78fb85fc5103c3fe66ffbe;
mem[496] = 144'h0105fe8a01980017008fffe4fe2dfff0fecc;
mem[497] = 144'h004e01eb00f7ffc6ffe1feedfe55ff8aff37;
mem[498] = 144'hfe6c0115ffac011a00f50120febbff0d001d;
mem[499] = 144'h009c0071feb00046ff13fe0f0120fef2ff16;
mem[500] = 144'h0151ffaafdb2ff41fdaeff97feccffc80070;
mem[501] = 144'hfedf0070017cfe6c0000019600b00076ff30;
mem[502] = 144'hfe7d0101ff5cff05fffefeabff490064ff2a;
mem[503] = 144'hfe69fe75ff0efe6a0148fe4e0147fe35ff3f;
mem[504] = 144'h009afdcc01c90243fe06ff11fe0900b3ffc8;
mem[505] = 144'h00f4ff98011cfff700c001d1fe0a0046001f;
mem[506] = 144'hff71feed02590012feca014dff910079fe5f;
mem[507] = 144'hfebafe01febd00abfeb6ff53013e0158fdba;
mem[508] = 144'h0109fe8ffde5ff8effe40133008a00c20105;
mem[509] = 144'h005f00ab0168ff56ff560073fef10143ff65;
mem[510] = 144'hfdf3006401a0ff63fed2fdbb012c00e2015b;
mem[511] = 144'hff4cfe97007afee3004fffbcffccfe9f0127;
mem[512] = 144'h00e8fbd8fa15026900ebfdee0584ff9afad2;
mem[513] = 144'h004efef8fc8ffe83fc20fba0019dfde9ffde;
mem[514] = 144'hffdc02710194ffe8f6bdfdb2fc5f018301e9;
mem[515] = 144'hfc82fa1bfd78025d0098ffca03a2ff8d009e;
mem[516] = 144'h0343fe08fca601650042fe1f017a0148fef2;
mem[517] = 144'h00cd0347fffe0054fd51fdf6ff0cff5800ae;
mem[518] = 144'h0171fce2fb3effe9ff2ffcb400e20034fd36;
mem[519] = 144'h037e011dfe0e01a30279fcc3016102c7fc45;
mem[520] = 144'h03cbfdcafb99fa13fae4fcea029cfe9bfd46;
mem[521] = 144'h03bf011ffdd9fe11fc95fa7601ea0284fdc8;
mem[522] = 144'h019c00d1ff99fffb016201d8fdcc0061fed6;
mem[523] = 144'h038afe6aff99019e022ffbbe008304c80097;
mem[524] = 144'hfa4dfc3b017fffe8fd89018306740167029c;
mem[525] = 144'hfd62f85ffe87051306f108f4fe08ffe8ff7a;
mem[526] = 144'h0137fc3efb66ffefff30fb8f0289fe86ff2b;
mem[527] = 144'h0190001cfc0ffe03fd02fc0703f90190fdd2;
mem[528] = 144'hffed0272060f02a003a203b80393fe86fd0b;
mem[529] = 144'h0152002e0636fe78fb0b008105fb0148fe8b;
mem[530] = 144'h011901ae0432fd91f400fcf4080d01af02ab;
mem[531] = 144'hf9aafd020657042a03c8026bfcb1fd4afd8a;
mem[532] = 144'h01e5012c0351002d0261029903f901c6fc75;
mem[533] = 144'hfddcff7f0097019dff43feac0317009effe3;
mem[534] = 144'hffd701cd059c0098fef5010f01bb0167fbb6;
mem[535] = 144'h02ccffc200a900fc039c008c02ab0216ffe3;
mem[536] = 144'hfd4901e606f7ff9dfd0b03c002ae0000fca3;
mem[537] = 144'h01590212029c0027001c034803a0003bfd73;
mem[538] = 144'hfd75fc75fd9d0389fd91fb6cfa86ff3e0216;
mem[539] = 144'hfdadfe3dffba03760554012a015100cdff59;
mem[540] = 144'hf436f6a1ffaf0226fce6024af60ef75cfd44;
mem[541] = 144'h07ff081f081eff5e027400220123043507a1;
mem[542] = 144'h00ccfec6089d0181fd8ffdd502fb0199fc2d;
mem[543] = 144'h018a0302052a006f0010027d02860273fe0c;
mem[544] = 144'hfe6dff6a0130fff6fdf0fe470050ff2c0114;
mem[545] = 144'h015afe56fdb4fe2a003c00860061fde8009f;
mem[546] = 144'hffea010bfe3dfe49fda0feb1011f00f1ff3d;
mem[547] = 144'h00c7ffa100f7fda8feb1ff16ff0bff51fe08;
mem[548] = 144'hff28fdccfe81ff46fe01002bffdbfdaa0070;
mem[549] = 144'hfe2201d3002f0072ffed004bfec901000057;
mem[550] = 144'hffcbfe1bff95fe17ffb6fe5700d8ff48fdb8;
mem[551] = 144'h0014ff28ffb1ff8a010e0134fe210113002e;
mem[552] = 144'hfee1ffefff4b00af0033ffe900c90022ff1b;
mem[553] = 144'h00eafdf4fec8ff8fff470032fde8fdde0127;
mem[554] = 144'hfec5fef2fe97fe270073fec4fe70fec8fdd9;
mem[555] = 144'hff9a00f0013b005400390138fddb0109feda;
mem[556] = 144'hffbdff770000009c0035fe740102ffb90056;
mem[557] = 144'hfe4500f8fef3feb8015700c2fe55fdebffa1;
mem[558] = 144'h00fafea5001a0104fda0fdf7ff640107ffbf;
mem[559] = 144'h0037fd9ffed3011afdf500dffec90034012b;
mem[560] = 144'h040302820141015cffbe02480391044201bd;
mem[561] = 144'h027d0236039900c4fefd0277fe38fd8bfa32;
mem[562] = 144'hfc04ff8802c8017fffb80437fac7fcf30062;
mem[563] = 144'h026dfb3dfd8effa1fcf70546ff69fea0fec5;
mem[564] = 144'h0619053a026101d5ff8afeb3033903f8018e;
mem[565] = 144'h0293012a020e02210019029601ca01d2012a;
mem[566] = 144'h0409015a0214012aff9b01040306ff07fb13;
mem[567] = 144'h05af02af031500b3ff41fd8a022602af00e3;
mem[568] = 144'h045e041b04dc002600e6ffffff37ff2dfd16;
mem[569] = 144'h060304f002c5008b002cffe701f8ff72fcde;
mem[570] = 144'hf6f0fbb901acff53fe8dfa8cfd5effd502db;
mem[571] = 144'hfe960232048901a90278f80d0211037103a7;
mem[572] = 144'hfa78f56eff4e01e900200509fa10fc330011;
mem[573] = 144'h02c2fb49fbc403d8009500f908c607560348;
mem[574] = 144'h05ec025f000002a1fdda01720180ffb1fb5b;
mem[575] = 144'h0471038c01dcffdeff4ffeb802ef017bffe4;
mem[576] = 144'h0505043402b103d8ff09ff4503ec06a60771;
mem[577] = 144'h021703f0fdab00c1feb5ff9e00c7ff8dfaa1;
mem[578] = 144'hfa73fc4b00a900c5feacfe1cf971f887fce2;
mem[579] = 144'h01620100fcb1021dfee5fe1702970a20028a;
mem[580] = 144'h0504063602d00215ff3500b0fdf8043104f6;
mem[581] = 144'h0020002401cbfea401f500defd49fcd40091;
mem[582] = 144'h014c01eb0012003afed6fce501cf0650fe1d;
mem[583] = 144'h006901480467ff6cffdaffe1014d031c0336;
mem[584] = 144'h03e0085302460100ffb1fdfa000500020034;
mem[585] = 144'h04fb079e054f001ffedbfd97005c03d30172;
mem[586] = 144'hf290fab20186fddefa1cfa5af792fe7303a2;
mem[587] = 144'hfe65026f0494fef6fcc1fd82fe7a027106b4;
mem[588] = 144'hfa7cfc64fed9ffa7fe1efeb3010b088efdf1;
mem[589] = 144'hfc6ef5e4f843036d03240126023201f8016e;
mem[590] = 144'h030101d2ff09007700c500c901260267fe46;
mem[591] = 144'h04c605de038c00380098fd1a000d0176043e;
mem[592] = 144'h011a00490217ffc3018dff48ff3a012f007c;
mem[593] = 144'h01950176fecb00950185feee00bbfecbff0d;
mem[594] = 144'h011dfe89010f002aff4c0042ffe3fdc0fea4;
mem[595] = 144'h0180fe1c00deff47fdf8ff3b0053ff0a017b;
mem[596] = 144'h013dfe50003fff30fefc0129ff5d0093fe97;
mem[597] = 144'hfee30118ff43fe77ff650072fef3fe7effac;
mem[598] = 144'h017dff8bfec600b5ff62004ffffa0118012a;
mem[599] = 144'hfe0ffe4dfe36ffc4fecafe190160ffaaff2c;
mem[600] = 144'h008d006cff29ff2d00ffff0a0123feca0145;
mem[601] = 144'hfebc008dfefffdef00ef004afe5c0123ff59;
mem[602] = 144'h006a0171fed8ff5301580042ffaa01c4fee1;
mem[603] = 144'h0222ff9cfea300060034fe410192febb00a8;
mem[604] = 144'hffa8fdcffe9bfdd5ff44fe62015dfedd00e5;
mem[605] = 144'h00d5feb501b4fe5bff4dff1b010cfe31ffc0;
mem[606] = 144'hfdcefe3501c6004d000dfdc2fe13011900c2;
mem[607] = 144'h00d4fef3fdd40078fe7bfeec014700f0ff97;
mem[608] = 144'hfd53000801acfc24fee80053fed8fdfcfe24;
mem[609] = 144'hff7402e406adfdd7fe6a001c00ae0298000a;
mem[610] = 144'h09d4094c07c6fe08ff7904ad086d059e0313;
mem[611] = 144'hfc5cfac300e8fedcfecd0204f9fdf470f799;
mem[612] = 144'h003f0041fed7fe50feea00dbff7efc87fcec;
mem[613] = 144'h0187007aff05ff1401020094fe3500a201c2;
mem[614] = 144'hff8e006a0153fcfffe970211fe84ff7afebf;
mem[615] = 144'h01ac00beff9effbaff6a012aff1afcbcfdcc;
mem[616] = 144'hff4bff7e02a0fcf4fe2b0157ff1700120036;
mem[617] = 144'hff92fdf000d1fc79fd20ff98fe4aff8bfe30;
mem[618] = 144'h0329fe7cff3104fbfe28ffb3034cfe61013f;
mem[619] = 144'hfedbfecbfc1e04eafdb9039d0128fcfdfec2;
mem[620] = 144'hfd9ff658fab1fea3015d01b0f6a1f88bfc0d;
mem[621] = 144'h0a900825088a02ef04ff048f070c06f507ac;
mem[622] = 144'hffc303510664fbd2fefa005e0112fe41ffe5;
mem[623] = 144'hfee0fef401ddfcda0025ff3c0087feb0fcd4;
mem[624] = 144'hff29ff3200eefee7ff82ff060100006200b4;
mem[625] = 144'hfdea0052005cfe95fdd1fdc3ff3afd840158;
mem[626] = 144'h0019ffc30143fee600a2fd0effe5016201f3;
mem[627] = 144'h00d9fe85fe7b0192ffbaffcd00f200330057;
mem[628] = 144'hff89ff9600bfff020005fecdfe710019ff38;
mem[629] = 144'h010f013c00930138ffaaffacfe8a0011fffc;
mem[630] = 144'hfd9aff34007e0195007201410169fe2fff80;
mem[631] = 144'h003bfef2008cff6401cdfef3ff1e005afed2;
mem[632] = 144'hff24fe260097fed1001aff2e014000f10142;
mem[633] = 144'hfeec00e100ebff42ff0afdb5fdc100e7ff19;
mem[634] = 144'hffc5fefa00e800c3ff63ffe2ff9affe10194;
mem[635] = 144'hffd8017c016fff68ff08feb3002aff84ff9f;
mem[636] = 144'h0007ffc2fe4c00c5fdccff400014fe83feb0;
mem[637] = 144'hff3fff53ff5dffe40035fe00fe87fd4801e3;
mem[638] = 144'hfd9dffa1013a01df00240100fe89fee00187;
mem[639] = 144'h009401f3ffe5fed3fe69fe86fe48ff56fed1;
mem[640] = 144'h04b0013c0139fc0ef7edfac003f8ff23fc8e;
mem[641] = 144'h0136ffa2fdd9f905fdd7048ffed2fdb6fdf5;
mem[642] = 144'hff38f99afdfe02b709530c02fb8f00690169;
mem[643] = 144'h02f40366005bfad4f979003b03d1ff86fe93;
mem[644] = 144'h01a104b40427ff1cf7bcf87cfedc00f9ffbf;
mem[645] = 144'h014aff75ff080129ff51ffa8ff13fef000bc;
mem[646] = 144'h028401d4ff16f7fefa3afd3c00ddfc0dfc03;
mem[647] = 144'h021d0174012a0189fb22fa1902e2ff52ff5f;
mem[648] = 144'h0300016800b6f8d5fd0bfd4afc68feb0fc5f;
mem[649] = 144'h04f304b1012ffa68fa7efbdbfeabfbf4fc26;
mem[650] = 144'hff1bfe8a0155006efcf4fc9700ba01d60251;
mem[651] = 144'h01d2012205270090f850f59000f901a900f3;
mem[652] = 144'h04b7097b03fef9befe0d03230347029401eb;
mem[653] = 144'hfc02f5eafc060a0d0a8305000675037003fb;
mem[654] = 144'h038ffee6fce5fa8dfbed003200b2fb2bfd80;
mem[655] = 144'h01aa04b80285fc0ff9edf97001c0fdc1fa6b;
mem[656] = 144'h000a00560070ffb6ffef017600000139009e;
mem[657] = 144'hfe4d013d017400c8011e0105ff0d0006ff6d;
mem[658] = 144'hff40009800d8fe5dffe6ffd00109fe2afe12;
mem[659] = 144'h00aa00c3fe9f00fd00dbfecdff92fde300f9;
mem[660] = 144'h0156fea4fe0effffffaafe2f013aff25ffd3;
mem[661] = 144'h0030005affd5009ffedc01bdfedb0037ffa8;
mem[662] = 144'h0138ff9300aefeb8fea2fe1bff2500ccfef7;
mem[663] = 144'h00ffff9bfe7bff5b0171ff2900bd00f80098;
mem[664] = 144'h00dcffd3fde9ff840150020200d5ffabff95;
mem[665] = 144'h0076fef9fe3bfe3c01360026ff0b008100c7;
mem[666] = 144'h0205feed018d0117ffa3ffb000ec0096ff58;
mem[667] = 144'h006bfee5001f00f30095ff34fe63fd96ffdd;
mem[668] = 144'hfde200d8ff60ffe2002efe07fffcfe75015d;
mem[669] = 144'hfef501d80146ff830064ff6efe2a006200b7;
mem[670] = 144'hfe3e006fff9f00b1fea8ff7500d60056ffe1;
mem[671] = 144'h007700db00b6fe00feca009700ab01f1ff44;
mem[672] = 144'h044602a2fe3cff4cfe43fd3a027a0266fba9;
mem[673] = 144'h063702eafd0b01800149ff98fdc4fe11fc34;
mem[674] = 144'h009cfcc1feb001150b010358f891015d0385;
mem[675] = 144'h00060268fe70fe1cffa0ffda02b9fcedfe45;
mem[676] = 144'h04650437016f019ffdf3fe85fd32042afe4e;
mem[677] = 144'h010700da00250013ff8a0191011c01d1fd56;
mem[678] = 144'h03020234fde700030192ffd0ff31009bfbad;
mem[679] = 144'h011d051b0228ff05017d035bfe320340ffbb;
mem[680] = 144'h04760178fbe1ff4e0304fd5801780132ff1a;
mem[681] = 144'h049a03ccfff0fedb0054fee4fcc2024bfbc6;
mem[682] = 144'hfa7b02b3ffe0ff4eff1402c1006001e700b8;
mem[683] = 144'h02630108037e005ff9e60232fddb0243ff3f;
mem[684] = 144'h030cfd6f0411fc870196feb60553fbb2ff82;
mem[685] = 144'hfd6cfd03fcb60334ff470635089d0144fef7;
mem[686] = 144'h01ad0493fe79fda80237ff81fe830058fd6a;
mem[687] = 144'h05880259fecdfe680045ffccffd10009fc6d;
mem[688] = 144'h025dfda0fc0efeddfed5fe6d015200fcfdb3;
mem[689] = 144'h00e1feb8fc9fffcffcca006e040c0100fd28;
mem[690] = 144'hfea702580107ffc8005d07fe0627ffe80065;
mem[691] = 144'h0160fb53f91a00d1fd2bff3a03ca041efe7b;
mem[692] = 144'h017200b0fd39fecbfe4ff991005d019b0331;
mem[693] = 144'hfc80fe26ff3afffb000dff94ff75fe58fccf;
mem[694] = 144'h00a3fc7af8c3fff7fd73fe4e047802d8fe3e;
mem[695] = 144'h022c0087fc87ff73ff16f938024104f30231;
mem[696] = 144'h021e0024fb010041fc7f022604d80236ff02;
mem[697] = 144'hfffbfff9fb0efeedfc6efa8f03060557021b;
mem[698] = 144'h0269ff8a0601fe0906c7fd1fff3100cf023d;
mem[699] = 144'h05e2013600ed01f504f2f5c700a5008b056c;
mem[700] = 144'hfb88fddefffc00a2fce10030038e034c019f;
mem[701] = 144'hffb2fc1ef9c902e5070dfe3ffc940069fbbb;
mem[702] = 144'h0148fd30f869feb5fc4dfe0a04d402d9fc9e;
mem[703] = 144'h009dfe95fbbb008efdf9fe78030304c8ff7f;
mem[704] = 144'hfee900a4fd82ff0e007ffe4cfd97ff3cfd86;
mem[705] = 144'hf9ee012dfe45002303e001b807220444fdd5;
mem[706] = 144'hfb73ff1efeb80022fda50442072bfcd6fd79;
mem[707] = 144'hfedfffccfee801bb036efdb90184028bfc86;
mem[708] = 144'hfdf5fe9fff14fe94fec20172ffc100e60272;
mem[709] = 144'hfd1bff50fc6efd70feddfdb8fbaafd22007e;
mem[710] = 144'hfd57ff6afebcff72038903ef020c05abfef8;
mem[711] = 144'hfeb5ff9bfcdafcedfe22fda5ff2101d00101;
mem[712] = 144'hfca7008effad01ad039c041905f501bf00c0;
mem[713] = 144'hfbb7fd02fd4f004c00f0025804260461ffbc;
mem[714] = 144'hff5d000aff93fcb100020038f87dfe2701fc;
mem[715] = 144'hfe210080fe09fed2fffbfe1afbc0fe5e0081;
mem[716] = 144'h007c012effac002201a9f8b90140fe93fe05;
mem[717] = 144'h0305fe05fe31fea4fd5ef8c1f638fe5afef0;
mem[718] = 144'hfae9ff07fe6cfff903870159054c03c5ff3a;
mem[719] = 144'hfd31ffddffc2000c006302eb016d01ebffb3;
mem[720] = 144'hff8101c107ab03ac00d8019e00b9003e015c;
mem[721] = 144'hff0a028e05bffd52faf9feb200faff77ff55;
mem[722] = 144'h05eeff260204fd65f868fc0202ec00d602b9;
mem[723] = 144'hff21feae02f202ff02fc023afbb200dd001c;
mem[724] = 144'hffdf017903ce00bc00b100fe0271fe50ff82;
mem[725] = 144'hff3402d2002b005cff7bfdfc010cfe560034;
mem[726] = 144'h00a9012c021efffd0038fee60005fda3003a;
mem[727] = 144'h01990133040b00fa048dfcbe020b0000fdbf;
mem[728] = 144'hffafff2d065efb7efb110111fed7fe7bfef2;
mem[729] = 144'h0140004304cd011ffd19fb94023aff10fe92;
mem[730] = 144'h02b7ff0c000f03b8fef9fdcb023501910228;
mem[731] = 144'hff68ff7c02c6030a016b02e1024d005bff4e;
mem[732] = 144'hfa9bfe10fe5eff0ffe4a02ebfac50140fe7c;
mem[733] = 144'h040e04c3051204b607a80899036203c508f3;
mem[734] = 144'h015d019a068ffeb1fcdafe9aff03fdd0ff2f;
mem[735] = 144'h018300b0042101a7fde1fe350113fe67fc50;
mem[736] = 144'hffe0feab00ccff3a00fc00230161ffa4003e;
mem[737] = 144'h011dfeeefea90038009cff9a0115ff9101c0;
mem[738] = 144'hfe2f00dc0038ff9f0082003ffedcfea8fe11;
mem[739] = 144'h01d0018c01dbfed6ffecffdefe5ffffe00fb;
mem[740] = 144'h0061fe40008dfe52ff83ff4efdeefe01002c;
mem[741] = 144'h019b015201dd0109016c0102014f00fa01bf;
mem[742] = 144'h010ffff5fe8601180049007dffceffe50145;
mem[743] = 144'h0102000800b7014901a7ffddffe601b3ff30;
mem[744] = 144'h006700ea015bff15ffc8ff69007efe11fe9c;
mem[745] = 144'h014600b301460043ffafff3f00cdfe160103;
mem[746] = 144'h01d60005ffe10107ff35fe8101bbfed3fdf6;
mem[747] = 144'hfe85fe85001000a700f900010069ff55fde4;
mem[748] = 144'hff7d009a0114fdc1fe76fe67fff50085ff9f;
mem[749] = 144'hff4300ebff07002dfe1fff230195ff5f004b;
mem[750] = 144'h007100130099010afe2901befea5ff45ff93;
mem[751] = 144'hff0b00af0026ff0efe67fee9fef3fdfafe47;
mem[752] = 144'h011c012e03f6fa1bfcc2ff5102d9fd6ffd5a;
mem[753] = 144'h00de00ae024ff855fab0010201c1ff96ff35;
mem[754] = 144'h0543ff46fe50fe3903ab0934014503bc01fa;
mem[755] = 144'hfdee04140511fb93fe4bfef90182ff72fdad;
mem[756] = 144'h00c201d6018afdc3fb21fbe0011ffef0fdf4;
mem[757] = 144'hfddaff5efef301c5ffd0fe9efe3dfe9fffe5;
mem[758] = 144'hfde9fff1009dfa3cfa8ffe5601d1fca1ffe2;
mem[759] = 144'h00ca005202dfff3bfcf5fda700bb0130fd24;
mem[760] = 144'h01c3ffb20234f861fc0c000a0134fc69fce8;
mem[761] = 144'hff2a01c40041f874fad3fd7a0135fd4ffc31;
mem[762] = 144'h052bfe0b01f4ffa1f997fc0300130166ff2c;
mem[763] = 144'h01a5ffcaffdd0148f6b3f959034000e7fe5a;
mem[764] = 144'h047d08000129fc42fc5b021dfd35fe19fc59;
mem[765] = 144'h007affe303ba06c10bc803f8021603390537;
mem[766] = 144'h001302bf0230f87cfa5cfd58024ffe1fff32;
mem[767] = 144'hff36006c0165f8a0fa0dfe13ffb8fd23fd1e;
mem[768] = 144'hff1f0152fb6dfe64fcc6fbd3ffc5009fff97;
mem[769] = 144'h008d0083fab5fe64feaffb56fc98ff5301ba;
mem[770] = 144'h0190fd12ff72034b072f02c9f98b00db0484;
mem[771] = 144'h02b001bffc1dfd83001bfa11059303d7ffb6;
mem[772] = 144'h027b002601b2ffa3fea8fdb0f984021d01eb;
mem[773] = 144'h00c70236fed4ffe200c2019dffe9fea1ffc5;
mem[774] = 144'h004f02bbfba8ff030054fba4fdc500e0ff51;
mem[775] = 144'hfee001e7008701effe53ffd3fcb3011e0169;
mem[776] = 144'h042cff6cfd4bfe4dff1ff9dffc95002902b5;
mem[777] = 144'h020a02da00befd82fcbcfb63f960ff8202b4;
mem[778] = 144'hff0a0110032600e6fe2906fd01ac029dfff7;
mem[779] = 144'h00830218fff5fedafaea035ffc63006f00c2;
mem[780] = 144'h04e506ce01bdfe59009afab50c0d08890441;
mem[781] = 144'hff65fa35fb4b055606ae09790105fe22fcb7;
mem[782] = 144'h01ec0127f961fd030097fb4cfe4cffd801f2;
mem[783] = 144'h00a20308fd6dfe66fdacf969fb57020b00f0;
mem[784] = 144'hfe3dfec2fd10fd5fff1e022a0013ffe4fbf9;
mem[785] = 144'hfc3a0029036dfed0fddd052a06e000caffb9;
mem[786] = 144'hffbc047c017201b1fbf006d609ad034f019c;
mem[787] = 144'h018bfd2201fbffb000a40108ff9d0065fed7;
mem[788] = 144'h0108fd59fddefdbdfd02009e05cf016d004d;
mem[789] = 144'hfd4bffe3fddafde8fdd5fe76fbfefe3fff90;
mem[790] = 144'h008dfc880041ff35fe37016403edffe6fd5a;
mem[791] = 144'hff10fcfaff97fef6ff6afb87055702e600cc;
mem[792] = 144'hfce100b800a6fc72ff29073f05a8fe95fca9;
mem[793] = 144'hfe79fdafff20fdcbfc7002aa0690001fff1b;
mem[794] = 144'h08ad0160039103330320fdbb02ab01dc00cb;
mem[795] = 144'h0277ff7affd502a30429fab7ff52003301f8;
mem[796] = 144'hfce5fe5aff75009f01c0038ef95ffa83ff9b;
mem[797] = 144'h0218022603a901630257f9a3fa3402fd02ab;
mem[798] = 144'h0011ff9cff96fe10fc74058a04c1018bfe11;
mem[799] = 144'hffaefc5bfda90053fe52029b03d40225fdc7;
mem[800] = 144'hff1ffe2300d0feceff7fff73fda7fef50104;
mem[801] = 144'h005c008afefefffdfd37fe79fe3cff9f00ef;
mem[802] = 144'hfff9ffe7fe4b00cd00fdffcafe830070fe0b;
mem[803] = 144'hfffb00710070fef30013fe5efd9afdf2fe0d;
mem[804] = 144'hfe2fff94fdf2fedb006a018e001300aefe68;
mem[805] = 144'h0116ffdd004affdbffcdff080073fe2301af;
mem[806] = 144'hff9afffdfe2fffacff57ff9400620022fff1;
mem[807] = 144'h007200b8fd3fff07fe99006afdfa013d0171;
mem[808] = 144'hfe69ff16003cffb900ccff290043ffb60000;
mem[809] = 144'h00ba00befef7fdd9fd800061003cfed7fd88;
mem[810] = 144'h0026febc008cfd45fe2efe0cffecfdcffe71;
mem[811] = 144'hffb6fdbafd57fde5003b00a8fff80025fddf;
mem[812] = 144'h0065fec0ff7cfda4ff7c005dfd6afdfaff13;
mem[813] = 144'hff86003300dafeb6ff17ffd0fdc9fe8dfeae;
mem[814] = 144'h00fb001cff90fe72fe4dfdc4fe510018fe87;
mem[815] = 144'hff38fd7bfd77fdb5fe24010affa6fef8ff44;
mem[816] = 144'h00befba8fa8f0117fd81fdb8055200ca00de;
mem[817] = 144'h02e8feb9fecefe7cfeddfdce0014028802c5;
mem[818] = 144'h0578028202190082031c02e7fe1f05f100fd;
mem[819] = 144'h0130feb8fda500e8fb22042f04b3fcaefe7e;
mem[820] = 144'h03c9fe7fff640178002efc78023b027401f9;
mem[821] = 144'h0211fff0ff17ff03001d00ddfe850093fe0e;
mem[822] = 144'h021a0052ff73fff7fea9005a002701ed0308;
mem[823] = 144'h031b0032fe0c019701810022023403ae0296;
mem[824] = 144'h03aafdaefd70ff74fcf5fbfe027802440146;
mem[825] = 144'h045c0001ff4a01fdfe2ffa31006404820094;
mem[826] = 144'h083201b5016b01030412018c002f00e5025a;
mem[827] = 144'h06880086011c0159034bfc44003500acff14;
mem[828] = 144'h0287fe8802b7fee1000403e30574f8d4005e;
mem[829] = 144'hfa03fe6dfcda033f02960746075f0259003a;
mem[830] = 144'h0201ffa0fe6500ebff5cffc2008effc0030c;
mem[831] = 144'h041500c9fd92ff9ffecefde1002a03a403d7;
mem[832] = 144'h002e0019017f057c050a042b011b04460690;
mem[833] = 144'h00e70034012506e2fecffd4802ca041b0506;
mem[834] = 144'hff1800880176007bf3c8f4e80277fcebffc8;
mem[835] = 144'hffc2ff6afe84081f03170598fe6f04c204f1;
mem[836] = 144'h006efeb4ff7e019b080504e5053900c9080c;
mem[837] = 144'hfd060000ffd4011bfffa00fafe93024b007f;
mem[838] = 144'h018e01ab019207300633005aff32038f05ae;
mem[839] = 144'h01e6ffcd014600030660026e008e01ab0327;
mem[840] = 144'h00080210fed8067dfe3100e30220041b0542;
mem[841] = 144'h013000edff6905d7031400a60323044307d0;
mem[842] = 144'hffd1fe1400d9ff76038f026c0060fc4900e8;
mem[843] = 144'h016cffd900d001dc096a041600f7fec402e7;
mem[844] = 144'hfb3afce0fe8c06e401a6009cffdf049f015b;
mem[845] = 144'h00a90002fc88faf8f855fbb0fb0cfdcffdca;
mem[846] = 144'hff2eff2ffded09240465fe5201b103600513;
mem[847] = 144'h016300b3ffb8084f0526025e023902e304c2;
mem[848] = 144'hfeabff8c03cc010100d1009bfb8ffcb6ff8b;
mem[849] = 144'h03ce026e07b100510168fce9fbe6ff2d0495;
mem[850] = 144'h0c0a03b1ffd4feee01a1faea0070065103a8;
mem[851] = 144'hfe70fd8b026e00f90338fff7fb39f79ffbcb;
mem[852] = 144'hfe15fcf50036015e0082034afd95fba6fdd2;
mem[853] = 144'h02b3033901d601e5015e0361046d039500a8;
mem[854] = 144'hffc9feb1067e020f02c3fca3f9a8fe230429;
mem[855] = 144'hfee3fd9301ab027202630330fe5cfad9ff75;
mem[856] = 144'h0161006b042d00cb0218f82bfcb1ff2302db;
mem[857] = 144'hff9cfd78019e00f200f6fda9f85afcb6012b;
mem[858] = 144'h00ff00cbfcb601a8fcb309b9052f01dcfcf3;
mem[859] = 144'hfc10fddcffad01570045088bff0ffb35fb1e;
mem[860] = 144'hff00f686fe6afef2ffcdfed90375f3f9004e;
mem[861] = 144'h07500c390a0f020b02b807da0b90041e04be;
mem[862] = 144'h01ca02d20811019a0244fe70fa31fdd8049c;
mem[863] = 144'hffb0feac02990338000afe6ff9d5ff4a0148;
mem[864] = 144'h030f03480028fe91fec9ff1cfab100030180;
mem[865] = 144'h0071032201560005029afd95f6b9fc940210;
mem[866] = 144'h00fe012402540531087c010af96cfa31ff0e;
mem[867] = 144'h028afe8e00dffca1ff72ffecfe5500b6048c;
mem[868] = 144'h025f0114043efe3cfc3c0072f9f9fa63ff1a;
mem[869] = 144'h0449001600de006803e502eb0080018dff95;
mem[870] = 144'h02f9ffde00a7fc46000000e7f998fcb80183;
mem[871] = 144'h01fefff0026efc58ff1c03d3fd90fdd70105;
mem[872] = 144'hff7e042d02e3fe750541fd0bf7aefe2800cb;
mem[873] = 144'h023600050455ff1e02dc013bf9c1f914ffd4;
mem[874] = 144'hfed701ec0133027afd300568097903b5fd0b;
mem[875] = 144'hfffd02a302c9fe20fade04260092fe27005f;
mem[876] = 144'h0319011200cffda00506fc9e0335023d07c2;
mem[877] = 144'h02bb0005fd5cfe41fd26054d067304d4ff2a;
mem[878] = 144'h00ac013a02effc8f0302ff6cfa11fceaff43;
mem[879] = 144'h025b029a0369fd1d012fff12f953fc7a014a;
mem[880] = 144'h033900e9fffef977f9fcfc49fd800143fde9;
mem[881] = 144'hff3fffb9fb1dfdb80062009cff5cfe95fb2d;
mem[882] = 144'hfadffcc1008802a90b700937ffaaf9c2fd98;
mem[883] = 144'h0240fedafe69f95cfbc1fa1403e0032efdff;
mem[884] = 144'h00dc00c00083ff08f841fcb0fa48fee1013c;
mem[885] = 144'hfe4dffa3013cffcd007a003cff2dfe91ffc4;
mem[886] = 144'hff13007afe6ff8a8fd05fd74fe1e0157fb52;
mem[887] = 144'hffdcff690251fe4ffb15fe8cfc5aff1a017c;
mem[888] = 144'hfe7e0087ff9cfb91026efd52fdfcfdf9fc28;
mem[889] = 144'hfd710240019bfc6cfd66fb61f9ab00c2fdae;
mem[890] = 144'hfb9a01a100bcfe3bfebb020bffea00560004;
mem[891] = 144'h002b02a40145fe52f81ffa1ffae7ff510080;
mem[892] = 144'hffbb027dfdbffc4bfebefb4004d706c000a4;
mem[893] = 144'h049cfe11fcee022c029402ce007b021800dc;
mem[894] = 144'hfeb300a4faf2fc52fd3afdddfdb9001bf956;
mem[895] = 144'h0063014fff61fa7afa80fe1afaee0090ff30;
mem[896] = 144'h01ab0287034c018001e90337030dff1f0205;
mem[897] = 144'h02a503f609cd0313fd90fa70ff0e00b5fbbc;
mem[898] = 144'h0419060a0607ff48fdc1faa50154ffbf00ba;
mem[899] = 144'hfcf1fcbc0121fef200d20251fb6efccbfe02;
mem[900] = 144'h04ff0160048a040b01dfff7c0118fde5fe71;
mem[901] = 144'h01e7011d04570053022cff45024b00ad010c;
mem[902] = 144'h039bff7c059800d502dbffacfc7dfe4bfdac;
mem[903] = 144'h031cffe9024bffe4045f02c0040b01effe1c;
mem[904] = 144'h013201d405bf0038fe20fb160140ff31fe96;
mem[905] = 144'h04f601e00704019cfe7bfc47feb70040fb9f;
mem[906] = 144'hfa61feeffddd02270434ff11039e0034ff80;
mem[907] = 144'hfe94fe51012c03a203e802b505a8fd79ff1b;
mem[908] = 144'hf963f22efc53014ffd6d0688fc0dfc29fde9;
mem[909] = 144'h0787090c0846ffbbfd1806350533049a083e;
mem[910] = 144'h0353014908440096fec2fe5afdd8ff8cfadc;
mem[911] = 144'h0485ffe6039c010502970056ff64fdfbffa0;
mem[912] = 144'hfd8dffbffef2fe98fe6ffe7a00530040006e;
mem[913] = 144'hff55fea8ff36ff7e00f4feaeff7bfee7fe1f;
mem[914] = 144'hfed5fe9affe3fda1fd94fee0fec7fe0e00e5;
mem[915] = 144'hffe5feb0ffe4ff64fef7fdfdff030059010b;
mem[916] = 144'h00cfff250075010f004e0079fe39fd81006c;
mem[917] = 144'h0057ff95ffe700a4ff9d0111ff1b014bffc5;
mem[918] = 144'hff52ff88ff88fdce0007fed7ff96ffbdfe8e;
mem[919] = 144'hff28001efe11ff8ffeebff07fd89ffde00d5;
mem[920] = 144'h0032feba005dffeaff5dfed0fed8ffbb008f;
mem[921] = 144'h010e0003feb3ffac009900c7ff5c0126fdef;
mem[922] = 144'hffee0097fff1feca01acfe2c00c2ffd90090;
mem[923] = 144'hfeebfdfb0088fd8b0108fd80ff6a001dff2a;
mem[924] = 144'h009600fefe74fdb7fe97ff07fe80ffe10043;
mem[925] = 144'hfd7bfd7fff0bfdb5feb5fda6ff68fe39ff50;
mem[926] = 144'h009b00a100b60038ffed0020ffb1fe5200d7;
mem[927] = 144'hfe880099012bfdb4ff4efda30023fec6ff47;
mem[928] = 144'hff7c03130125034e046f041601f904b10556;
mem[929] = 144'hfd520188ff41019e010efb370361035afee1;
mem[930] = 144'hf8fdff92fe19fdb8f4c4f95501e3f9f20048;
mem[931] = 144'hfd5501a7010a055f05c8fe79fef509c4030f;
mem[932] = 144'hffe500ab00500289043e0436ffb300c407a9;
mem[933] = 144'h000efe87fe94fff3fd71fdd8005000b80297;
mem[934] = 144'hfd2a00b1020a041804cefebf026f06e70434;
mem[935] = 144'hfeaa011400f1ff0704ab01fe001000c502fc;
mem[936] = 144'hfd9202ee014601b8ffb400b403a3050b066d;
mem[937] = 144'hfff9041c03d3024805390345ff8706ae0703;
mem[938] = 144'hf729ff9200c3fd38fd7901b5f47ffed702f8;
mem[939] = 144'hfd04fee302cefdde002304d7fd1001b405fb;
mem[940] = 144'hfe430300fd600085001efcb3033a0a1cfe18;
mem[941] = 144'hff88fbd9fd76fd4b0137fdfbf82afe58ffd3;
mem[942] = 144'hfce80244013702fe01c4fe79fef4072403d0;
mem[943] = 144'hfe55034100eb036b0465ff5b0243064a052f;
mem[944] = 144'h00ca0051fe1aff3c00b0fd6c009fff7dfec0;
mem[945] = 144'hfd9bff1f009bfe3cfe8efe57fdddfe980042;
mem[946] = 144'h0041ff9fffaafdebfeef00cb0118ffb8001b;
mem[947] = 144'hfebb0097ffad00e6ff80008afd8efeeffde0;
mem[948] = 144'h00edfdc0002b001300e8fe0bff8c00d1ff90;
mem[949] = 144'hff82008f002d00f900b301c1ffd501270073;
mem[950] = 144'hff6f005ffd7efdccffaefdf7fd7fff320014;
mem[951] = 144'hfd76fdf7fecffed50012fea0ffbcff42ffbe;
mem[952] = 144'hffabfe7dfde3ff740020fd6cfda6ff5afed9;
mem[953] = 144'h0121fdaefefdff4cfdc3fe46fdde012000d9;
mem[954] = 144'h00f7fec900e6febafd89ffc100940059ff8d;
mem[955] = 144'hfdd700f7feff00580106fdb8012f0060fdec;
mem[956] = 144'h0139ff60ff4ffe0fff1dffacffc2fe40feca;
mem[957] = 144'hfe57fe7bfe2dfed6fe530079ff6f00b6fe20;
mem[958] = 144'h00cffe53ffa9fee30085ff44008300c2ffde;
mem[959] = 144'hfe21feb1ffb2fe40ff85ff2dffcafec8febc;
mem[960] = 144'h0045fe64ff3f0174008fff6c0023fdeafffe;
mem[961] = 144'h0161ffd30140010bff3b00bfffb5ff4e0016;
mem[962] = 144'h002dfe620120ff7cff4f012bfe51ff8afe35;
mem[963] = 144'h00b7000301b000a0fe200168013c00630039;
mem[964] = 144'hfe8600fbfdccfe99fe16013000f9fe5bfee3;
mem[965] = 144'hfeb201d9018bfebe0066ff0e0165ffecffee;
mem[966] = 144'h013200520036fec8feb3fe3d016eff9aff56;
mem[967] = 144'h00e1feaafe2dfe7bff5101a5013900310173;
mem[968] = 144'h00200158fe70008cfe07febbfef0fdfdfe3c;
mem[969] = 144'h00a9ff76fe6c000b0068013afee4fdc6015c;
mem[970] = 144'h005000c6ff6a002bfe8a002f00dd0113011e;
mem[971] = 144'h0066fe00fde200f10025ff45ffcb0052ffad;
mem[972] = 144'hfe9a0072ff00fe6600f201040178010dfe31;
mem[973] = 144'hff04fdeefe0c00d9ff93000aff9e0120fe76;
mem[974] = 144'hfeb7005c00d80039ff1700b1ff5001340100;
mem[975] = 144'h00d4ff59fdc5014200ad017fff9cfef30020;
mem[976] = 144'hfe52fd64fd66ffe8fd00fd7afe3bff190012;
mem[977] = 144'h0004fd51fddafe45fd34feb0feec00a4fdce;
mem[978] = 144'hff820182fdceffa1ffd6fd8901500047ff97;
mem[979] = 144'hfe20ff19fedc0058fd51fe8100fdff53fe3e;
mem[980] = 144'hfd1cfffcfd6b00e2fff4fce9ff5afffbfcdc;
mem[981] = 144'h0153ffc60147016fff2d019bffedfe41fe8e;
mem[982] = 144'hfd30ff85ff2a00dbfd58000efd00ffbdfe14;
mem[983] = 144'hffacfde1fd31011efe8cfe66fdd6fdd00079;
mem[984] = 144'hff53fdd2fdbd00fdfee80048fd51ffb1011d;
mem[985] = 144'hfeb1fea6fe7d011f0000fd6fff3301ab007d;
mem[986] = 144'h01e9ff0bff2d004efe0f01010043fe0f0055;
mem[987] = 144'h01e7fe21ff62fd91002b0299fe63fdf2fd0e;
mem[988] = 144'hfcb0006bffb2ff16fd87ff7b01860024fd78;
mem[989] = 144'h001afef0fd1a0040fd63fe16ffdffd5c0007;
mem[990] = 144'hfcf4fd3cfdd0ff8ffd26fe83fe19015fff15;
mem[991] = 144'hfdb8fe7dfe0b012efce10041fe5900d800df;
mem[992] = 144'hfe24fd4ffc4cfda8fd35fe8d0290fd7afaec;
mem[993] = 144'hffc8fe5ff917fd7702a4058b03d3fe2afe92;
mem[994] = 144'h02930164ffae040d0a1d09a2003604c60128;
mem[995] = 144'h03a704fd02c3fba6fec300dc05190015fddb;
mem[996] = 144'hfecfff71fc9bfca0fa77fe45ff22029cfc64;
mem[997] = 144'hfd4cfe06fdc3fcf0feadfe90fd9dfedcfecd;
mem[998] = 144'hfeb40168fd43fdf8fe8402fe046afdc70040;
mem[999] = 144'hfd5a00e4fd6b001afb5bfc0700c30277fdc8;
mem[1000] = 144'hff13fdb5f791fe67024003a2034cfe77fcf0;
mem[1001] = 144'hfe43fdb2f9aefd44fce1024701f2ffd7fcb4;
mem[1002] = 144'h08d903900133ffba04c700f101e5046800c0;
mem[1003] = 144'h063303860156ffa3fd5cf8a801210157feeb;
mem[1004] = 144'h0d1c0dd30502ff6c0099004b03dbfe400243;
mem[1005] = 144'hfa1ffa0c00a600fd00e9fb86fa1afeb6fa8e;
mem[1006] = 144'h00b5ff85fc61fe3100c602de01d2fd49fedd;
mem[1007] = 144'hff7dfea1fad7fd79fbbbff9f02e0017efed0;
mem[1008] = 144'h03540033fe75ff5502aa009cfdb200e6fbc3;
mem[1009] = 144'h007dfe56007101a90035fc5d017e0206fd2c;
mem[1010] = 144'hfe070106015d0049fdb4001905c1051d036c;
mem[1011] = 144'hfe7afabefff6013c0122fe0dff8bf967f95b;
mem[1012] = 144'h032b0103fe00ff0801450154fd5c0287fafa;
mem[1013] = 144'h017300b1ff19fdbe004dff150152034cffcb;
mem[1014] = 144'hfea7fe25fea2ff6e0111fdabffb6025ff9e4;
mem[1015] = 144'h0281ff15fff5fe8101500164fc6400f5fd66;
mem[1016] = 144'hfda9fed1fd25fff9ff28fe9fff91031dfb97;
mem[1017] = 144'h01a9fd6dffa9ffb9fefcfcc9fed1010bfc4a;
mem[1018] = 144'hfb7e0380012b019704ba0455ff0c01f2ff04;
mem[1019] = 144'hfdccff83015f0161042a0197fda901effe1f;
mem[1020] = 144'hf4d1f13dfca80310ffa8ff7f0129f912fea5;
mem[1021] = 144'h0ce309be07f0fdddfd1502880274fc33ffdd;
mem[1022] = 144'h0144fdf0fd65017c0210fcfc002d046dfc32;
mem[1023] = 144'hffaaff1fffb0018b009efee6febe011efbb9;
end

always @ (posedge clk) begin
	q_a <= mem[addr_a];
end

always @ (posedge clk) begin
	q_b <= mem[addr_b];
end

endmodule