`timescale 1ns/1ns

module wt_fc1_mem6 #(parameter ADDR_WIDTH = 11, DATA_WIDTH = 144, DEPTH = 1024) (
input wire clk,
input wire [ADDR_WIDTH-1:0] addr_a, 
input wire [ADDR_WIDTH-1:0] addr_b, 
output reg [DATA_WIDTH-1:0] q_a,
output reg [DATA_WIDTH-1:0] q_b
);

reg [DATA_WIDTH-1:0] mem [0:DEPTH-1];

initial begin
mem[0] = 144'h02f103be021d023b008d02d900db035202fe;
mem[1] = 144'hfe6702c0046afef90000ff3a02d6016bfe19;
mem[2] = 144'hfd39fde0ff0bfc8bff40ff86fdf5f7c3fac3;
mem[3] = 144'h022f0543003fff09004c0478013c03bcfeba;
mem[4] = 144'h010003ce01d302d7ffbdfff200ca0281029a;
mem[5] = 144'hfe4bfe2b0083fd00fce1ff490081ffb4fd28;
mem[6] = 144'h0242057c039302f2025d01a3020b01dcfde2;
mem[7] = 144'hfec8005803f001fbff11017ffd3b020600be;
mem[8] = 144'h010c065203af00640162011800a7ffe1000b;
mem[9] = 144'h02d8050f050f03070135fe8c01e9ffac01d3;
mem[10] = 144'hff94fb30f8e8fcb700b50134ff5dfd29005c;
mem[11] = 144'h0051027dfffd01b7ff48006203220122044b;
mem[12] = 144'h00fd0644fc05faf4ff55fefc008d0528fec8;
mem[13] = 144'hfb9ff93ffafc00d0031401a4fbeefc47018a;
mem[14] = 144'h004404a2037efe83022400fa017bffa8fce9;
mem[15] = 144'h007103c6040800c20161ff7b003f041f01a7;
mem[16] = 144'hffd6013cfe8efe03ff96012f005bfef1feae;
mem[17] = 144'hfe4601d70150ff0cfe8c00ca00090034015b;
mem[18] = 144'h0003ff7fff8e01a3ff1d006aff01019f0129;
mem[19] = 144'h012100edff790224ff7901d4ff2c0067ff61;
mem[20] = 144'h0067ff2dfee5fec7ff7600fe0018002e00c4;
mem[21] = 144'hfe26007afe9afe42006f0152ff41014f01a9;
mem[22] = 144'h00a3ff41015fff30ffb4018d0143fe5fff99;
mem[23] = 144'h008d0170fe80012dfe86ff7cfe810219ff35;
mem[24] = 144'hfec9ff5efe8dffbefe74fdeb00bbfe7dffef;
mem[25] = 144'hfefa00d900690136ffabff0e0063ff4aff67;
mem[26] = 144'h00b8ff3d023901dd0244fe1c001f00f500b9;
mem[27] = 144'hff49fee9fe1c00d3fe2aff05febaff7cff50;
mem[28] = 144'hffe3feac016cfe34ff8a002fffd3fde500a4;
mem[29] = 144'h005bfeebfe3d0067fdf101c8000d00c9ffa2;
mem[30] = 144'hffca00e300e1ff70000b01e2ff8101070214;
mem[31] = 144'h0030fe0901fd0087fe8affef0179fde7009b;
mem[32] = 144'h0121fe55ffe3007dff23fecbff290022ff76;
mem[33] = 144'h01610193ff1dff94010a008300e4014c002e;
mem[34] = 144'h001001930052feedfed3ffddffedfe81015e;
mem[35] = 144'h00f1fece00ccff0ffe31ff8d01950058ffd3;
mem[36] = 144'hfe5cff78fe67fe790181fe9dff3e011afe58;
mem[37] = 144'h0031ff9001deffa8fe53010100d0ff6300e1;
mem[38] = 144'h003a00a8fe32011afee7015efea0ff1eff53;
mem[39] = 144'h000efe6dfefa01c2ff3101720185fee60114;
mem[40] = 144'hff90fe9cff31fe29ffcf0089fe18fe650173;
mem[41] = 144'h01c0ff4b0070ffd200bdfe590119ff1400f3;
mem[42] = 144'h00eefe95fee3ff9b011b004c0139fe66ff05;
mem[43] = 144'hfea1fe82ff4b00d1fe37003f013201090051;
mem[44] = 144'hfdfa002fffbcfedbfe14fddafe39ff2bfed1;
mem[45] = 144'hff600025fef9fe9a0155fea3fe8900b60083;
mem[46] = 144'hffd8ff41fe970176006fff54fe9301d6ff01;
mem[47] = 144'hff2dfe38ffe6ffa1015b00feff3cfe450184;
mem[48] = 144'hff15fdd20083ffeaff7dff19fe94fdb7fd81;
mem[49] = 144'hfe3cfe3afdee007a0015fd72fd8bfdb5feeb;
mem[50] = 144'h0055008300f3fed7febe0060fe65fdacfe1b;
mem[51] = 144'hff64fe8200b0ffb4fff7ff760015ffe2fd73;
mem[52] = 144'hff42008700c5fde20079fde3fe6f0076fe31;
mem[53] = 144'h015c00c9014d00ae000d01720158fed50046;
mem[54] = 144'h00b9ffe2fd8bfd59003efea3fd5900fdff25;
mem[55] = 144'hffdefe70fea70047fee8ffa2005a00c9fed0;
mem[56] = 144'hfe6dfe44fefc00e5ffc5ff80000bfdf700b1;
mem[57] = 144'hfdf6fe4f004aff4cffdffe06fee5009cfdb2;
mem[58] = 144'hfe5a00c5001afe15fffffe510027ff91ff31;
mem[59] = 144'h00eaff17ff21ff96fd93ffb7ffaffdf9fe31;
mem[60] = 144'hfe58001bfef1fd6b00f8fe3dff3bfea0fd61;
mem[61] = 144'h00fffd63fd72ff01fef2fe69002bfe58fefe;
mem[62] = 144'hfe150053fe5eff36fe1b009afe8a0003fe46;
mem[63] = 144'h00210025fdf4fedb005e00f4fdb8fe110091;
mem[64] = 144'h04ba04ba0139014c00a401ad012a0175fe23;
mem[65] = 144'h008f00acfe5e00d1fc84fe5bfde9fa52fb7d;
mem[66] = 144'hfc78fb13ff86fee4f975fe7afa9bf8defeb8;
mem[67] = 144'h03c3002afb0a01d0016701470197fe9b00fb;
mem[68] = 144'h023f03aa0391fd4800830057fbb7ff74fda1;
mem[69] = 144'hfe12013f0000021cfd23004d00a80057fe45;
mem[70] = 144'h051701affc91000fff690140fea0fde0fe70;
mem[71] = 144'hff8704670298ff1301feff97fe1800a4ffcb;
mem[72] = 144'h038e01040029fe58fb400175fd2bfc66fc2c;
mem[73] = 144'h039d040bfe44fff2fc45fd74fdc1fce7fb5a;
mem[74] = 144'hfe93fabffffbfd9000fd0062ff9304f40768;
mem[75] = 144'hfe7c00780497ff0401cdff8b009903390161;
mem[76] = 144'h03cd0011ffca0558fe79ff2f02d2fed90032;
mem[77] = 144'hfe14007300cdfd8905a30503004900cf01cc;
mem[78] = 144'h021a02b6fba2008400ec001bfe5afdadfd11;
mem[79] = 144'h01cb03feff40ff43006bff2dfef50059ff2d;
mem[80] = 144'h00a0fedbff4301040023fe4a01bcfecefef5;
mem[81] = 144'h00c8ffd500c2008d01bfffabff05ff7affc7;
mem[82] = 144'h00ceffbefe6900ce00630035ffc1ff55016d;
mem[83] = 144'hff56ffa90120ffa3fefa00cc00af0049fe2d;
mem[84] = 144'hfeb7fffc01a3000e005a00cafdd100c5ffcb;
mem[85] = 144'h004bfe78ff9d00dffe5200bdff5ffe3600b2;
mem[86] = 144'hff7bfe8a004000d6018dfe23006d0117ff41;
mem[87] = 144'h0181fe84fe720004ff0400b900faff310025;
mem[88] = 144'h0076006a0189ff080023009200d6015aff3d;
mem[89] = 144'hfff00186ffc4ffc3ff83ff12fe6bfebeff2a;
mem[90] = 144'hfe5dfdd60108ffb0ffc9023ffe210007011e;
mem[91] = 144'h020500f2fe77016b00f301fffe37fe48ff7b;
mem[92] = 144'h00a0ffe4ffd7ff660083fee9004bfe3aff6f;
mem[93] = 144'h0002014efe2400c1ff73004d0179ff4fff3e;
mem[94] = 144'hff090137fe93ff3e004000350152ffecffd2;
mem[95] = 144'hff720206ffa60062ff6b010a009ffef5ff5f;
mem[96] = 144'h011404650150fc8fff2d036904c4063b0343;
mem[97] = 144'h03fd057eff59001b019a01da046204000304;
mem[98] = 144'h04100456fcc7067400a90125fe3cfc99ff11;
mem[99] = 144'h039a043f00f2fa82016503290438050dff1c;
mem[100] = 144'hfe68011f035e01c3fc15ffaf0062051a03e5;
mem[101] = 144'h00d6010902e5ff7704a9015802cc02e802a1;
mem[102] = 144'h03bb0406052afc74feef033c03e20499025a;
mem[103] = 144'hfc17016d03c5fdd3fe0b015b017703b102ea;
mem[104] = 144'h04c205ec01dcffc9ff08029b029d02260242;
mem[105] = 144'h02a1046e03f8009001710328047702be063c;
mem[106] = 144'hfed2fb2f00f10581fedfffaffd5cfef70121;
mem[107] = 144'hff8efb360546013bfe52007ffcce01810620;
mem[108] = 144'h02f504e202ccfe4500ab026601b401ecfc1b;
mem[109] = 144'hfd87f9abfd4dfb5bfc280031fe73fd66fe37;
mem[110] = 144'h04a1037a01cafcf8010702c2054b038d0188;
mem[111] = 144'h040303de031000cafe6101de032504b0035e;
mem[112] = 144'hfebf01f7fe8bfe56010b01e200f9ff1dfed4;
mem[113] = 144'h00cdfe44ffa2ff06ff9c00b400520060ff41;
mem[114] = 144'h0188fe7dff310085fe37fecd0087013e00bc;
mem[115] = 144'hfe2d0031fe34022e0185ff5a0242ffbafe6c;
mem[116] = 144'h0036fe55fe14fe50fdc0021eff56ff6800c8;
mem[117] = 144'h013101060161ff2cfefc002900ffff75017f;
mem[118] = 144'h013201e000d8fec8015afeea004a00270127;
mem[119] = 144'h00400061ff7701a800cdff68ff92ff1c000f;
mem[120] = 144'h01fd0063ff0501faffdcffc800ebffb5fdde;
mem[121] = 144'h0071ff34fe2afde700220113fe1dfdfafebd;
mem[122] = 144'hfe7cfebefe61ff8cfedbfdf6011cfee6fddb;
mem[123] = 144'hffcf011dff3dfeeb0168ff5a012100bdfec6;
mem[124] = 144'hfe6bfde001470148ffcbffb2fe4bfede00d3;
mem[125] = 144'hff2f00b1ff2d015400060242016300f50069;
mem[126] = 144'hff7a013c0058fe81000100d7fe5bff10feba;
mem[127] = 144'h0102ffc6013f0050ffd6ff5600e4fefd0073;
mem[128] = 144'hff7700550011018901db0040fdc4fd79fd56;
mem[129] = 144'hfe8aff50014a00030212ff6dfdf600fd003a;
mem[130] = 144'hff04050701a4fc3e0175004f02fe003dfc50;
mem[131] = 144'h0029feb2003b01d8fd9cfcb3fcd400360191;
mem[132] = 144'hff8700a2fe3cfe8401bc01c4fe30fe05fe91;
mem[133] = 144'h01f400cafe06ffa900d5fe39ffc101dafffa;
mem[134] = 144'hfe11ff59ff8c0325ff48fd3efecbffdffe9b;
mem[135] = 144'h028bff7bfeb9ff8f00c00102ff27fe80fdf5;
mem[136] = 144'hfd43ffa5ffc0ffaf03cdff56fcf3fdaffef5;
mem[137] = 144'hfc99fe7dfd6b000901d20123fddafeddfd41;
mem[138] = 144'hfea0020905dcfa73ff570129010604320162;
mem[139] = 144'hfe7c01f201f2fcc600740283ff770081fecf;
mem[140] = 144'hfeebffb701b00279ff1affb1fe36014f036e;
mem[141] = 144'h08be0815fe9b00ee03d200a802a90291fdfb;
mem[142] = 144'hffbfff8d01bf02b20111fbd6fba5ffdaffe1;
mem[143] = 144'hffe2ffcafdbeff090387fe96fd8dfd05fce6;
mem[144] = 144'h01090025fde1fd8c0054ff240455fe74fb7e;
mem[145] = 144'h0094fd34fb94ffa8038503bf0442008c01cc;
mem[146] = 144'h00f6ff7601a404450019063a014e0827072c;
mem[147] = 144'hff1a018dfb5900f60298ffb8ff7bfb36fc17;
mem[148] = 144'h043e0053ff7efd6d0317ff26058b0269ff8e;
mem[149] = 144'hffb5007a028d01a101dbffcf001b033002e3;
mem[150] = 144'h011f008ffbdffe3804d504bb040efdfdff14;
mem[151] = 144'h015d000f00fbfb0b0221ffdf01aafebbfe84;
mem[152] = 144'h0432fd8afe45001f028304ce06da033302ee;
mem[153] = 144'h040cfd4afdedfdc60227040f04b0006dfeea;
mem[154] = 144'h01f1026406a6fda3013a0106ffc80193fb49;
mem[155] = 144'h00d400e20183fa4d005800adff5701c9f8ca;
mem[156] = 144'hfd1affc2f8fc072601acfe29fdedfdbdfbfe;
mem[157] = 144'h00e60650043efc46fe2e000c016300d801af;
mem[158] = 144'h0138fda0fbbbffb7060d034903e2fda2ff2b;
mem[159] = 144'h0228ffe3fe73ffd8033b0145050002440197;
mem[160] = 144'h010f0221fd3601ae03050018fdd4fbe20031;
mem[161] = 144'h011500d3fbfd06eefd7afd4afbd9fc030030;
mem[162] = 144'hffe5fb0d0bbc0460fad40134ff2e047e0522;
mem[163] = 144'h03fd0237fc3c080d0260fb53fc80fe89fdc5;
mem[164] = 144'h0306017b0468fccd05cd0285fec1fc880085;
mem[165] = 144'h008d01cc00f600d602c7018c00ab00970220;
mem[166] = 144'h014b0302fc38025c0418ff95fe8efbb7fdae;
mem[167] = 144'hff8403a3fd97fcc402c4027ffec5fc23ff75;
mem[168] = 144'h0179ff20ff730362ff5f0094fac7fd6affc8;
mem[169] = 144'hff680168fe66021305c2021afdc9fc79fd80;
mem[170] = 144'hffc8fe5e0918fe1e00ec02e002e0ff66fb0a;
mem[171] = 144'hffc1fff10540f9d5049204a50254fb2bfc83;
mem[172] = 144'h00bcfff4fbf40bac006802c4fff1fe5201ab;
mem[173] = 144'h0198054705e0ff970452fcf0045a08ba085f;
mem[174] = 144'h02a7fff1fe0a026f01a6fe4afd50fc44fefd;
mem[175] = 144'h02df01fcfcdfffc603a301c3ff48fad7fe8e;
mem[176] = 144'h016effabfe72ff2cffea00900103fe86ff29;
mem[177] = 144'h0064000a013a0006fff9004dfff1fef800e0;
mem[178] = 144'hff2affd200b7fe2cff39fe520167fe81ffb6;
mem[179] = 144'h00ff014cff6202190235ff5fffbd00b5ffba;
mem[180] = 144'hffa2ffd1fdd3fdc800cb00b4fe1c0075010c;
mem[181] = 144'h018e008900cb0149fe5ffe5d00c3ff260114;
mem[182] = 144'h00aafe41fe3cfe9affce020eff3bfde3fe42;
mem[183] = 144'hfea8fe32fe2fff11009e0096007c0052fed6;
mem[184] = 144'h01ea000bff5600d2fe53fee8020701b7000f;
mem[185] = 144'hfecffea4fffe0107fde600e700daff6cffd2;
mem[186] = 144'hfdf7fea700a700a7fefdfee9ff51006a001b;
mem[187] = 144'hff390141fed5ff40fe3200acff07feabfe05;
mem[188] = 144'hfe4bfe37fe03fe5affdafeb8ffdffe7cfe85;
mem[189] = 144'h012afeb4ffe4ff17014b002efff7ffa800ff;
mem[190] = 144'h0012fe4e00b4009fff9bfef9009001c7fed3;
mem[191] = 144'hfed6febe00f4ff7a00d0fe7c023500b50116;
mem[192] = 144'hfe73ff5f03ed01ec018401fbfe25009b02cc;
mem[193] = 144'h01e40489048a035600ffffc50079ffbfff57;
mem[194] = 144'h021f01f7fc73fc2803c0fe28fe82fc4ff79c;
mem[195] = 144'h01d200660211ff75f9b6ffff00200252043f;
mem[196] = 144'hfdca00e4011b03de02d0013ffeae00fdffe1;
mem[197] = 144'h00c7ff4c00a3fd1cfef0fee7007d00fd0072;
mem[198] = 144'hfee40130043104ec002100c501d1ff5a0288;
mem[199] = 144'hff4bff98ffe4018a00810104fe4201d80008;
mem[200] = 144'h023901c203c9044f00930229fffffe24fe38;
mem[201] = 144'h0210024f023502e402bc0140fdc3ffe7ffcb;
mem[202] = 144'hff95fd40f973f9c4ffa4ff77014d04bc01c3;
mem[203] = 144'hff49fe46ff7d009f0284ff0400cc059a0094;
mem[204] = 144'h0295011e04def7eaf95afd30ffa2ffd50148;
mem[205] = 144'h00040021fe4a004a01f101250015fd53fcc8;
mem[206] = 144'h013700ab04c904f6fe44021c01d60193fffa;
mem[207] = 144'h00f0ffe9025e04570007fee90008002b01f5;
mem[208] = 144'h026f0092003702c4ffd0ffbcf86afcadfdc6;
mem[209] = 144'hfd80fd830217044ffdf9ff69fd66fc7bfc40;
mem[210] = 144'hfd3000a90528fe49fd62ffbb03b80596ff67;
mem[211] = 144'h0006fd50ff0105a0fefafe08fc68fa2a0172;
mem[212] = 144'h01be0371fe3201af02fe00b9fdb9fc0ffb98;
mem[213] = 144'hfea5007600bcffe0fc9eff8dfe39fe9aff9a;
mem[214] = 144'hff9afe0ffdcf0492fe19fc9dfa88fd9bfe04;
mem[215] = 144'h024201a0fc01055000d8fef2fe96fd6dfd41;
mem[216] = 144'hfaeefe0bff9cff0fff46feb8fa60fa15fb64;
mem[217] = 144'hff8bfe89fdc300effe90fd3bfb3ef98ef855;
mem[218] = 144'h023804ea0261039f0330026300c6085705e1;
mem[219] = 144'h02ad04c0ffaf025e0252001c02200118fd3f;
mem[220] = 144'h0125ff960294042c01cfffbcfe70fe7506ae;
mem[221] = 144'h02960474020104ea041f0158012b059d0429;
mem[222] = 144'hff33fd4800a503d0008cfe54fac1fe17fc9b;
mem[223] = 144'h02bcff0dfce602a40136fe13fb45fa82fc3b;
mem[224] = 144'hff4aff5cfd930034ffb1fde604760235ffb4;
mem[225] = 144'h0095ff83ff0dfed0ff1a006f01d5ff73ff93;
mem[226] = 144'h00cb031b02470066ff3b02edfe3dfe2c0441;
mem[227] = 144'hfdc2ffc6fea5fe7bfee0fd190359fd91fe3a;
mem[228] = 144'hff9cfe380083fc5dfe53fc99001b026eff43;
mem[229] = 144'hff9fffc40205feb5fea301590010026d0227;
mem[230] = 144'h0018fe46ff41fede005afd660378013eff1e;
mem[231] = 144'hfdd600ba0020fd80fe85fca4025d0220ffe8;
mem[232] = 144'h039f018efd0500c0fea2fe87045402d80031;
mem[233] = 144'hffc80072fe4afefc001efccb05eb0274ff2d;
mem[234] = 144'h0303fab7fed301810475ff4cfec5fe4efd97;
mem[235] = 144'hfe6cfb8afdd0007c0190f9b8ff1001bcff3d;
mem[236] = 144'hffae0271fd7d01f1fbc501650081004ffbbf;
mem[237] = 144'hfb68fe4000f8fe210081fd6ffb8cfc9aff35;
mem[238] = 144'h01b0fe71fef1fdfc0166ffe103d8ffa5ffc2;
mem[239] = 144'h00c80009010dff90ff0dfe96029302b0fed3;
mem[240] = 144'h02ac0348fe4cfe7501150400ff24009a000b;
mem[241] = 144'hffae00a8faddfe5700a4fa9a00680100049c;
mem[242] = 144'hfb7cf927ffa3036dfaabf9d2ff31004706b1;
mem[243] = 144'h0407026dfefb0137038302df0216029dfccc;
mem[244] = 144'hfe0d025d022bfb18fe66003a007f00cd031c;
mem[245] = 144'h00ce022f02f1006902f6ffc0010101c500a2;
mem[246] = 144'h0145018efc2dfc4e0289ff8a00c9fe08013f;
mem[247] = 144'hfe5801ba03f4fcb700cb013cff3f01df017a;
mem[248] = 144'h000e034bfd23016600aefcddfdd40201057d;
mem[249] = 144'h011101f4ff32fd00034002bffbfafe890532;
mem[250] = 144'h029201f9089f03ea013e02210175fc1b0138;
mem[251] = 144'h02b006030824fdac017d01d40083fbac01e8;
mem[252] = 144'h02f400affd40066105330552002d011bfee2;
mem[253] = 144'h004afed401cffd33fb98fecb03780662fec8;
mem[254] = 144'h021800abfba4fc0e0270fd8b0125fe9eff94;
mem[255] = 144'h027a033400eaff1b013a0134ff7dff3801fe;
mem[256] = 144'hfd37ff3a0227ff25020bfede01f101caff41;
mem[257] = 144'hff91ff8afda0fe770513fe7e0454044e0480;
mem[258] = 144'h02500235faf902e20453fec80351018005f8;
mem[259] = 144'hfd4500d102b5fa03fc34fff2025701fbfec7;
mem[260] = 144'h01b4fd0cfec800f8ffb3fff206c901ce0362;
mem[261] = 144'h00b80096ffae00ae033b02fc029e00c8fff8;
mem[262] = 144'hfd40002d0255fb2c00d5ff96010c012f0344;
mem[263] = 144'hfcd2fd36ff0a0042ffb8003a042bff7300f7;
mem[264] = 144'hfe8e003dff39019203d8fe7e061d0389051f;
mem[265] = 144'hfeb6fed2fddcfdf304e3005a045a057f0532;
mem[266] = 144'hffc5fc69fd08fc9bfe86ff20fefcf5eaf906;
mem[267] = 144'h01eefd09fb4fff6e00f600bc0083faf8fb6a;
mem[268] = 144'h005500effbdbfb8c00b4012400d3fd7dfe50;
mem[269] = 144'h0497026d05170386faaaf91e053703f8006f;
mem[270] = 144'hffb2fe250039fdaa0080fda9025201ae0330;
mem[271] = 144'hffbafdf201bbfe0ffff301ca010a021300ca;
mem[272] = 144'hfff0031e0152fd6c018f037d02120569070e;
mem[273] = 144'h031e02bc00cafff200e8fcf5ffdb0117011e;
mem[274] = 144'h020400ed042b0846fc79fe12fc1efa5f034d;
mem[275] = 144'h030e02cffd49fdff0364040404690492ff0b;
mem[276] = 144'hfe450444035efd14fbf80232fed603da054e;
mem[277] = 144'h018a008a00e4027b02f60248014b01ab00bc;
mem[278] = 144'hffb905690007fdfc036202d80237029e01ac;
mem[279] = 144'hfd8a00e60515fdf1fe8dffe5fed4020405e4;
mem[280] = 144'h033a069c0101013f01d301f00048035a0374;
mem[281] = 144'h009802a305640171025300fd01ff02680722;
mem[282] = 144'hfdf9fdeb04340182fd59fef2fda6f8e2fc84;
mem[283] = 144'hff0bfd7a0586fc95fd7c02effe82fc7606a9;
mem[284] = 144'h03d2042cfe4b012c04c7024201cc0501fb2e;
mem[285] = 144'hfd39f96cfdf7f9d0f9b7010800850572054a;
mem[286] = 144'h01d501ec01f7009f00c401a901b3005d0069;
mem[287] = 144'hff5104a802f1ffba00100410003704d704cd;
mem[288] = 144'h012afdf702eb03b80145fabb00ceffcffd69;
mem[289] = 144'h0159ff2dfd79fc56fcebfef103b80003ff40;
mem[290] = 144'h02d9ffacf8edfd47018003bd02b107cc0682;
mem[291] = 144'hfee0fc6e02a6fdc6fb30f87602ccfdd6fc43;
mem[292] = 144'h025bff20fe5e01cf008efc7103fb02e5fdcf;
mem[293] = 144'hffea01c9001501ee023dff11ffb701400181;
mem[294] = 144'h00b5fe34013cff07fd70fb4a0089ff98fdc1;
mem[295] = 144'hfe48fe8600f40277fff8fe2b014501e2fbaa;
mem[296] = 144'h0036fb53fb87ff0901faffea05770175fd24;
mem[297] = 144'hff73fe3bffb400baff59fe01028402aefcd3;
mem[298] = 144'hff7bf63df658025a02e90216fcdbfb7affc6;
mem[299] = 144'h0094f96dfd0e04800460fd79ff4dfdc0faf9;
mem[300] = 144'hff82fb7eff69fc8bfd810259027efba3fff8;
mem[301] = 144'h03f104cb0f2b08a6015dfb0c040d02aa0524;
mem[302] = 144'hff8bfdbbfd55fd7ffe0bfbf002a9011c0007;
mem[303] = 144'hfe6bfdf90137ffe7ff94fcdd01f60189fcf4;
mem[304] = 144'hfea300270023fe20ffd0fed4011dff3b006f;
mem[305] = 144'hfe87fe78002efe8201580122ffdd015e015f;
mem[306] = 144'h0096019bfde5008affb4ff45feb7fef0ffbf;
mem[307] = 144'hfea6fdf7003f0146fef7004b01780087ff5c;
mem[308] = 144'h014b011a0120ffacfe430109ffb000f3ffea;
mem[309] = 144'h01b70162ff0300efffdc007dfed701c500c1;
mem[310] = 144'h00d3011ffe1d0122ff33fec6009cfe94ff0e;
mem[311] = 144'h00180118fef8004100b2ffdfff18ff4bfedb;
mem[312] = 144'hff980026ff50ff2900ecfebe000000a20082;
mem[313] = 144'h01b4fddbff0bfd9800b9ff6f001e00b5ff16;
mem[314] = 144'hfdc0027801bbff8efeb6fe7ffe7dff5f00b3;
mem[315] = 144'h00cd019fff20fe7affbfff6bfddf01b3005c;
mem[316] = 144'hffcfff21008bfe69ff1100faff9a0018ffb3;
mem[317] = 144'h00bbffd30040fdf90059fec4017900e400fb;
mem[318] = 144'h000dfec80043fe5a00feffe8fe2efe62ffca;
mem[319] = 144'hff64ff800043006cfe64006e00f3009ffdc9;
mem[320] = 144'h028e0530005600bf01d701bffe63fb77fff6;
mem[321] = 144'h010dfdfbfcd101080119fb27fba0fc9d008d;
mem[322] = 144'hfb4df95a00330255fc91fe29005400bb04cd;
mem[323] = 144'h030d04bafcc10313049c0211fe82ffb300cd;
mem[324] = 144'hffdc02ee02d4ff65026e0190ff91fb72ff90;
mem[325] = 144'h0093027fffe900a9ffccfed3fe1300f6002a;
mem[326] = 144'h00fe0278fabd005504e6fd4dfe2dfe04fd37;
mem[327] = 144'h040105080038fede03c803a6fec7fda9fd06;
mem[328] = 144'hfe04ff86fff90074ff4ffe40fa1ffe4e00b4;
mem[329] = 144'hfee000ddfec7000803080103fb5bfbdbff94;
mem[330] = 144'hff34046703fd029e0105029f020e0351fd91;
mem[331] = 144'h033805b105d8ffce03dc040c04cdfd4ffee3;
mem[332] = 144'hff9f016200fe072e050801a6ff0e019203e8;
mem[333] = 144'hff87ff25032801270046ffe402aa05710004;
mem[334] = 144'h013bff1efaae031a02b2fe33fc20fe5e0084;
mem[335] = 144'h03a2018bff63018f03a501effdb3faeafe64;
mem[336] = 144'h0054015b021401c00142ff77fb21ff73ff24;
mem[337] = 144'h0158017f01be04df017a000bff00fe040026;
mem[338] = 144'h02ac0258011ffea700aeff0d01550035fcb8;
mem[339] = 144'h0187fe6d03f90272fce7fdd10078fda003ef;
mem[340] = 144'hfeb3fdddff2f00fe028203c6fe3cfc75fd08;
mem[341] = 144'h01ceffd801cb02400151ffd0fff400c40073;
mem[342] = 144'hfee100aefe930158fe43ff0cfbd3ffc4ff71;
mem[343] = 144'h02ff025bfda6022400d603fb001afdbefdd0;
mem[344] = 144'hfdefffb6002100c502fa006cfb5bfe8a00ad;
mem[345] = 144'hfecafed7ff9b00e200a40093fa6dfbc9fe63;
mem[346] = 144'hff8000040021fb67fdb702f000b501d201ac;
mem[347] = 144'h0020ffecff4cfed3001e01770250fefefe06;
mem[348] = 144'hfea4fdcb036dffd9fdc5fe7aff1301690499;
mem[349] = 144'h058003cd019c004903b4ff7803f60269fe5f;
mem[350] = 144'hfd510162ffa40485ff86fe12fc3fffae0144;
mem[351] = 144'h002c0079fff6018802320123fe1bfd1cffd6;
mem[352] = 144'h0245043901a9ff63ff110120043b01130115;
mem[353] = 144'h04f8021a01cb03c902e10569fee30048fff8;
mem[354] = 144'h05b90240fea803ee02d8034afd460298fc3b;
mem[355] = 144'h030e0198fd0eff4900ad00d40317fd3dffcd;
mem[356] = 144'h0053025a022cff6e01310041003a0241026a;
mem[357] = 144'hfe1bfcf501d60120fd51fdf3ff3f002dfefa;
mem[358] = 144'h0484049d0170033c014405d9021d0173feb9;
mem[359] = 144'h017301360105010dff45ff4a032f014a0070;
mem[360] = 144'h05f50346029b0359022606000089031cfe6d;
mem[361] = 144'h0777047d02da02af021b04a9027001eb00cb;
mem[362] = 144'hfefefc6301bd00dfff0300c9fe2b05f10384;
mem[363] = 144'hff13fe7501d5fffffe590093febf0503026e;
mem[364] = 144'h02fcff64007000fefda1011d0319fee50092;
mem[365] = 144'hfa9f029cffc7fc1ffdee006f040a00f102c4;
mem[366] = 144'h04a402edff49047301d3064602bf013300b0;
mem[367] = 144'h051404e1011e01e301a1050802dc01e3ffa4;
mem[368] = 144'h0119ffa7ff0300b0fe7400f9ff65ff240025;
mem[369] = 144'hffd4feaa01ba015601df013101a20107007a;
mem[370] = 144'h0142003eff9700aaff110012feb200c801c6;
mem[371] = 144'hfdcb017afffcfffbffad00f60170ff400038;
mem[372] = 144'h00e7feeaff40ff0cfe790018001ffe9f0123;
mem[373] = 144'h014dfec7feedff47ff83019d00a0011a011c;
mem[374] = 144'hffadfffafee6fe38ffed015d01b1ff24febc;
mem[375] = 144'h016b010f0176ffb1ffd9fe96ff5c000900a9;
mem[376] = 144'hffb2feb4ffd101a3005901de01c4fecdfeac;
mem[377] = 144'hfeaafe6eff70008900af00720038fe2cffbe;
mem[378] = 144'h007d0019ffa4000901a40013015cff1cff92;
mem[379] = 144'h008b010c0043ff9ffef50021fea3fe39fe10;
mem[380] = 144'hfebfffbeff37fdeaff2afecd00bbfeacfeb3;
mem[381] = 144'h0040fff300f3ff2d0107ff8b0105ffab0059;
mem[382] = 144'h0167005ffe8c016ffe64018200e9fe1f015c;
mem[383] = 144'h00570184fdf20180003f0011004bff1f0083;
mem[384] = 144'h035fff79feddfd60ffedfdabffbf0057fea3;
mem[385] = 144'hfd90fd55fcd6fdd7feb1fd65ffc3fcfafcf1;
mem[386] = 144'hfd90ff46fedeffdb00a4ff62fda9fdfafeab;
mem[387] = 144'h0111fd8b002efef700d000c7fe28fffefffc;
mem[388] = 144'hfe9401a2fda0fdaffea1001bfd9e0063fde7;
mem[389] = 144'h0038ff65fe83fef2ffd1ff13fe58feb4ff48;
mem[390] = 144'h009a004ffdd4fd3f00b9fe11fed6fe67febb;
mem[391] = 144'h02c50160ffa90018fe08fddafef1fe64feb5;
mem[392] = 144'h005dfd040054003dfe8d005cfe6bfe9cfdd2;
mem[393] = 144'h00b4fd5bfcd70075007f0059fd3afe32fcec;
mem[394] = 144'hfd8a010801dbfe35ff59fe67fee3013affc4;
mem[395] = 144'hff5a0014feaafd6fff0ffdd0fe2b01e20082;
mem[396] = 144'hfe48fdd8ffa8fffc010efe02ffb0fd4afe98;
mem[397] = 144'h0099fed60039ff6dfe4fffd3fd4ffd35001a;
mem[398] = 144'hfe40ffc6fceffe84fe67ff1dfd32ffd6fd54;
mem[399] = 144'hff9e0045fd760005fe9dffbcfd28fd77fd6e;
mem[400] = 144'h034f01fdfee101c2ff00fd6b017bfe9bfd1e;
mem[401] = 144'h02bd0088007703acfdfa03d5fdd3fdcffd5e;
mem[402] = 144'h0284000004ce0083001e03ecfd88060afd34;
mem[403] = 144'h02510078ff41061bfdf500b000a8fc34fe8c;
mem[404] = 144'h027303ec002c00a70339003f015a0033fc0b;
mem[405] = 144'hfcacfcd60035ff38fc3cfdea00f2fd7d001f;
mem[406] = 144'h05ea01c4fde00443ff5a01c80045fbfffd03;
mem[407] = 144'h04bd04c7ff67009a02780129016d0311ff92;
mem[408] = 144'h0351fe0701070039002a03b9fba6fc09fc46;
mem[409] = 144'h0568036e017701f3038e0281fe55fc1bfc7a;
mem[410] = 144'hffbdffffffb0fe1dffbcffba0025049d037c;
mem[411] = 144'h021e00f100b0fdd40364fdfbfeca0298fdab;
mem[412] = 144'h02f6fd68015605f5fbab0021ff11fed0031b;
mem[413] = 144'h000104d000b8fccd02ee0053059d09730622;
mem[414] = 144'h0210007800c8038a01ef012dff02fefeff0e;
mem[415] = 144'h0579035ffd8702bf01cb02170107fe07fd27;
mem[416] = 144'hfbf9ff8cff0bfe6ffdd2fe13fb3afea4fd6a;
mem[417] = 144'hff4a0031ff01fbcffce3ff9bfdfafe3bfe0f;
mem[418] = 144'hfc69fdeeff2bfbb1ff2efdc2fe85ff030195;
mem[419] = 144'hff71fcb7fd95fcd4006bfe71fdcaffcefdd6;
mem[420] = 144'hfd36fd95fbe7fe02fcb4fcfafc9cfe1bffdb;
mem[421] = 144'h01760038fe38019bff79fefb013efe3cff65;
mem[422] = 144'hfeaefdbafe50fddcfe09ff1cfae8fe5ffef8;
mem[423] = 144'hfebcfc5a0050ff9dff17fce9fc4afc60fdc5;
mem[424] = 144'hfedeff4ffd2bfcdbfc06fd1ffc95fe11fea4;
mem[425] = 144'hfe98fdf5fef6fd5cfca4fd33fcc6fec2fcde;
mem[426] = 144'hfe68fc77fcff0028ffcefcd0fedbfb10017c;
mem[427] = 144'hffb8fc2ffc26fd9f00bcfe60ffdef9ebffb0;
mem[428] = 144'hfdb5feb2fdbcfcb101b8fe89fd0cfe1cff16;
mem[429] = 144'hff45fe8a00db00490131fe8fffb10063fe3e;
mem[430] = 144'hfdbffd20ff7cfad2fc60ff10fde5feeb0058;
mem[431] = 144'hfd20fccafc49fe73fdc6fe1dfcd0ff2afc85;
mem[432] = 144'hffe5fecd0215013cfee9004900790023ffa7;
mem[433] = 144'hff6dff21fef1fe54017501d6ffcbfe4aff3a;
mem[434] = 144'hfdfdfdfe00c600530045ff79012a014f00c3;
mem[435] = 144'h0081febcfddafed2fdd5014afebeffda0153;
mem[436] = 144'h0139fe3afe2dffaefe3a010aff470046011d;
mem[437] = 144'hfeb2fffafe360029fe5200160177ff41013b;
mem[438] = 144'hfdfafeab01cdfeb80074006400dbfdc8ffc5;
mem[439] = 144'h003d0060013501c901730063fedd00e401d2;
mem[440] = 144'h00170037fe0afe7f007400a50179013a0126;
mem[441] = 144'hff7a00fa011a01850065001bfefd01420093;
mem[442] = 144'h0033017ffdee002dfe20ffec0081ffc4ffa0;
mem[443] = 144'h00b2ff29ff9300f0002e009e0077005ffe01;
mem[444] = 144'hff80ff79005a010cfeb8fe8d00f000690156;
mem[445] = 144'hffbffde001750120fe9afe2000abff8e01e2;
mem[446] = 144'h01cbff3c0093002effbf018fff650211feef;
mem[447] = 144'hfe32ff6f023afda5ffed0032ff79fe10ff53;
mem[448] = 144'h002bfee8ffbcfedbff03fff4fdc30129febd;
mem[449] = 144'h006e005c017cffe5015cfff4006a00b701b4;
mem[450] = 144'hff46fe1bfdcffe36ff56001100b4fdf8fe8c;
mem[451] = 144'h00c1011501e8009600d8ff9c00ad00fdfddc;
mem[452] = 144'h009bfffeff94fe07fe6f017d01750106fee8;
mem[453] = 144'h01ce00a2011201b8ff230123fe98ff51ffd0;
mem[454] = 144'hfe7afeb0fef200be00fa01420154fe48ffc1;
mem[455] = 144'hff0800da016e009afff6ff8500b3fe4ffe55;
mem[456] = 144'h015a00990098ff2b0153ff9900c300030128;
mem[457] = 144'h01450053ff42ff59003eff4d01bbfe430007;
mem[458] = 144'h0003ff87fecf013b008300c8008ffe6d0105;
mem[459] = 144'h0107fe37fe95004600db015a00010147fffb;
mem[460] = 144'hff72fe41fdd7fea20127fe18017700c6ff60;
mem[461] = 144'h010f009dff83ffc9fe73010cfef6013bfe6b;
mem[462] = 144'h01a8ff02feddfe830048ff2d0177ff4dfe09;
mem[463] = 144'hfe94ffef014e014ffe3bffa3fe13ff30fe0f;
mem[464] = 144'hfac8fcb302a802b401bb01b2febb02ba0327;
mem[465] = 144'hfe9905f3089c02bbfe36026afff00086fda1;
mem[466] = 144'h02b005af055dfb38010f0185ff78f880f72f;
mem[467] = 144'hfc39ff7602f6040cfa7000a7fe7d04c003e7;
mem[468] = 144'hfca8fd6d005e00ad007aff71fdddfe41015f;
mem[469] = 144'hfefbfdb6fd3bfe6c008b0101ff57ffcffe08;
mem[470] = 144'hfc41029204000586001902f6fea00398025c;
mem[471] = 144'hfc93fdd8fec1039a0138fe2cfddf005c0300;
mem[472] = 144'hfdb0041206ee0296010203f9fe69fe49fed4;
mem[473] = 144'hff7e02fb0478031fff640110ff2fff5600c1;
mem[474] = 144'hfeedf99efa0dfade003800b10361fea0ffc1;
mem[475] = 144'h0142fb80feb000b5010a0013002d0355049a;
mem[476] = 144'h007404df0632facff83afda2fe3c049b02da;
mem[477] = 144'hfafdfcb1f86cfb6d05be04fffc56faae0072;
mem[478] = 144'hfcb9026b046a02eefeda0042ff0602bcfe63;
mem[479] = 144'hfcb201e30277030bff0c01cdfd100357039b;
mem[480] = 144'hf8b4fc06050b01fbfcdbfe70f9a201e803f0;
mem[481] = 144'hfc84039807f3fc87ff460418fee60254fd95;
mem[482] = 144'hfd0c0728fefcfa2a044d023f008bfa04f5b4;
mem[483] = 144'hf7dafec304aafec6fd6c03c1fbf407bf0449;
mem[484] = 144'hfb97fdbb00aa0335fbd9ff0cf97ffd0e0124;
mem[485] = 144'hfe520045fd33fefbfd41fe70006dfcceffae;
mem[486] = 144'hfa9efda1057b0014fd3a04f3fb5905020331;
mem[487] = 144'hfde2fb8d014602f7ff46fd82fb92010f0328;
mem[488] = 144'hfa6f045d0775fd3eff9e0295fe27ff54fc6d;
mem[489] = 144'hf8a5005306c10202fa74001cfd8a019cfe73;
mem[490] = 144'h021cfc8efc100479ffa5fec6020805290d81;
mem[491] = 144'h013ffa7bfefc04a8ff3efb9101a203a708ff;
mem[492] = 144'hfdf008fe0419f505fd7cfed701af086a04de;
mem[493] = 144'hfe9bfca0f73d060c037e0470f740f5c5fef0;
mem[494] = 144'hf7c4011c06ea0242fe5204f2fd7c022c006b;
mem[495] = 144'hfc30ffb105a702dffb550157fc820291002c;
mem[496] = 144'h008dfef300e8ff8601340070ffa80150fe9b;
mem[497] = 144'h003b01e8ff6c0085ffb5ffe5ffb1ffd4fe47;
mem[498] = 144'hfe2e00aa017a0184ffb6012c01b0015b005d;
mem[499] = 144'h0124feb40027fdcfff03fef50110014dfe05;
mem[500] = 144'h0242ff30ff5900ce00a1fe4701bdfe7a005d;
mem[501] = 144'hfec9feb2fe8dff93ff20fe5dff3d01d7fe89;
mem[502] = 144'hff73010600470000ff28012d0160013ffe74;
mem[503] = 144'hff6c004cfe61fe9cfe33003a0129006ffe8c;
mem[504] = 144'hff0d0023fe020117ff60ffe7fde4ffe3fe7d;
mem[505] = 144'hfe2f00f000dbffdcfdaffe57ffc7ffb7000f;
mem[506] = 144'h0081fea6ff8a0050ff7afe2aff97fe91ffc1;
mem[507] = 144'hfe59fddd004eff97ffdcfe63fdb9fff8011b;
mem[508] = 144'h010500a00016002dff880003fec2fde9fec1;
mem[509] = 144'h0099ff1601adfecdff87ffa5003301a80151;
mem[510] = 144'h0139fdd6fed0fea300b80161ffd3004400ec;
mem[511] = 144'h01b001550085ffa1fe760123ff9aff3d0069;
mem[512] = 144'hfa0cfac800510030ffacfd2ff919fed00395;
mem[513] = 144'hfb4dfe3106a50094fd2d0509fbdb00a3fd3f;
mem[514] = 144'hfe4d06410644f813029804ce0024fd96f68f;
mem[515] = 144'hfc1efd7c06d70297ff520159f78b04160400;
mem[516] = 144'hffe4fbe1fe4c02750104fd38fe17fb2b0151;
mem[517] = 144'hfcfeff1cfdbbffbffe37012d00a8fecafee6;
mem[518] = 144'hf858fadc04d8019bfe2e002cf99d0110010b;
mem[519] = 144'h0061fd1bfd3a0272fe8bffc6fe32fdfd00da;
mem[520] = 144'hf90f0050053c00b7ffa20113f82cfeb0fd7f;
mem[521] = 144'hf908fe3e012602e3fe3dfde1fa41fe3f01a3;
mem[522] = 144'h01f00201fc9a01a10244009102c20096071f;
mem[523] = 144'h0333fcfbfbe905100312feae0432ff3d0688;
mem[524] = 144'hfbf50345079cfffcfb33ff45fe2a06f2ff83;
mem[525] = 144'h0237fd90f89802e1029d01bdfd88fc580000;
mem[526] = 144'hf94afdae050b03a8fea3ff47f969ff6001aa;
mem[527] = 144'hfa02fd1d005803b6fd0a002ffc30fda503d5;
mem[528] = 144'hfd41fb1c0028012cfeddfc75fe15012fff5d;
mem[529] = 144'hfd01fc5c01b7fbdefdab02ee03e603ddfe23;
mem[530] = 144'h038505a1fdabfd07024e04650655049e0040;
mem[531] = 144'hfbfbfc72043bff91ff0bfbbeff44fd1bfcce;
mem[532] = 144'h017bfe51fd0103640257fb9e01c802d1fd0e;
mem[533] = 144'h0043ffeeffb0006900c9feef00e701240001;
mem[534] = 144'hfd06fdd00010fd62fd03fafbff30013c0084;
mem[535] = 144'h014efbebfd7a02a9013efd67ff9bff85fe1d;
mem[536] = 144'hfdb8fcfdffa1fee5fd1a00110135010aff2d;
mem[537] = 144'hfea5fd69fdfcfe6bfeeafd16036802f8fc65;
mem[538] = 144'h0117fc67f8e5063206b7014eff08fc590485;
mem[539] = 144'h02aefaf0f8db041b03e2ffb20107fe6f0002;
mem[540] = 144'hfeedfc15011efe1f00e0033f0132fc3aff1e;
mem[541] = 144'h0766044b052c088d0109fba4029a0461062a;
mem[542] = 144'hfd39fd0100a6fc97fd05fc84010803130120;
mem[543] = 144'hfc47fc71008b003dfde0fe6eff6cffeffc74;
mem[544] = 144'hfe7d005f008300ddff13ff57fe13fea0014b;
mem[545] = 144'hfd9ffe0efe74fee8fecdfe160143ff1cfe65;
mem[546] = 144'h0070ff39fe13ff2300c2ff880054ff06000a;
mem[547] = 144'hff70fff5fdf1fdc4ff6ffed70035ff56fedc;
mem[548] = 144'hfe29ffb3fe43008c012afdfafe50fdf5fecb;
mem[549] = 144'hfe53fec300ccfef8ff57001601b7ff62016d;
mem[550] = 144'h0077ffba004700dbffe2fe00fdd1feacff6d;
mem[551] = 144'hffbefdfffdf6ffeafe34010e009bfec7fe47;
mem[552] = 144'h0101fdbd0062fe410095fe05fe130146ff4f;
mem[553] = 144'h0077003cfdf2fd9bffd900adfedfff03015c;
mem[554] = 144'hffea0043ffd70001fe9900c9fecd0085014e;
mem[555] = 144'h006900e1fe8bfe3e006200cb0136002d0028;
mem[556] = 144'hff190098fe13002400a7ff4e00f8fffafea8;
mem[557] = 144'h0106fe16ff2d010cff96007200b9fe0afe9a;
mem[558] = 144'hffbdfe15fed4feaf00b2fe84fda3fe45fdc3;
mem[559] = 144'h0066ffd0004a013e0085fe6000dbfe22fea1;
mem[560] = 144'h002ffe2ffe30fff902a4ffd504e5fd4cfcb8;
mem[561] = 144'hfe2ffddff9fcff410212ff040453027a0224;
mem[562] = 144'h000ffd71fc3b02310014017302340455067b;
mem[563] = 144'hff57fed6fd08fc9400bafe09fe61fe34f8d3;
mem[564] = 144'h00d4ffacfceefb7d01c1fe200206021ffd55;
mem[565] = 144'h010a02e60095029bfe980230ff8300f2ffe0;
mem[566] = 144'hff2cfc74fadffc6c02a2fe65023afdd6fd73;
mem[567] = 144'hfeb6ff1c00dcfb910061fe5300b1fecafc78;
mem[568] = 144'hff37fa43fa14fe3e0378ffd404d304e40016;
mem[569] = 144'h006efef5fbd2fad80153fe6506710338ff03;
mem[570] = 144'hffbcfe9f0133fd1500f5007cfdb7fbbafb49;
mem[571] = 144'h012d0234fed9fdc9031cfde3fda7fce4f95e;
mem[572] = 144'hfeb2ff1ff5bb013a0448fef3feb7fc70fd10;
mem[573] = 144'hfe9804fb05bf03d1fc47febc006e03e30072;
mem[574] = 144'hff9efe0ffdc0fb13040ffef501e0017fff46;
mem[575] = 144'h0274fd03fd57fb36ff42001a037300e6fd59;
mem[576] = 144'h01a201daffcfff8101d9ff93039e0030fe25;
mem[577] = 144'hfff400befe47010501e4ff5702e3ff61fd76;
mem[578] = 144'hffd4ffb9fd43fcb7003e028afcb5fb350213;
mem[579] = 144'hfe8c005cff92ff930224fd0b028e013dfc58;
mem[580] = 144'h00aa023e0169feaf010d0065011901bcff0e;
mem[581] = 144'hfed50086ff59ffe1fe92fed2fe78ff18feba;
mem[582] = 144'h030201af004effa8016801d102a5ff67fee2;
mem[583] = 144'hfe0502970017fcb8ffab012bfe4ffe70feac;
mem[584] = 144'h013dffddfce2febf022d00df006801fa00dc;
mem[585] = 144'h02580324fd53fd0401c5feea02210144fed5;
mem[586] = 144'h00cdfe790122f9ed00d8ff81010ffe3f0102;
mem[587] = 144'hfcb4ff270009fbb7038aff720099020ffe4b;
mem[588] = 144'h011a036bfc2c0093fcf0fd16ff33fe4dfb95;
mem[589] = 144'hfef700520066fcc90274045cfefcfc0afb0d;
mem[590] = 144'h003f0270fce6fea803dd00f300d6fe30fdcf;
mem[591] = 144'hff0801a1fd7efe260081fed6031b02c9fe6a;
mem[592] = 144'hfe5aff79fdd900b9ff3f0179ff2b008dff54;
mem[593] = 144'h019f00b5feb9fecaff9300e70165fff9fe62;
mem[594] = 144'hfefcfe35ff83feddfea7fdfb0189fe8bff3f;
mem[595] = 144'h01630052fe72fe33ff3e00d000d2fe980078;
mem[596] = 144'h019101d001dc002afef0feb5feeefec8013d;
mem[597] = 144'h00e700fb0168ff1300bcfe4e0013fe5cff20;
mem[598] = 144'h011dfe8500b50036fedcff0cfff3ffd50061;
mem[599] = 144'h00e0fff3ff40fed9ff9fff0efe2e001f0075;
mem[600] = 144'h014e0082ff22ff920068fe2d0038fdc9ff35;
mem[601] = 144'hfdc5fe0200f00113001f00e7fe67016200db;
mem[602] = 144'hfdc40022febd0132015efe7affaeffde01ef;
mem[603] = 144'h0151febf01f5feeb0149014100c7012bfffa;
mem[604] = 144'hfe1cfe740168008efdb800c90135fe3dff11;
mem[605] = 144'hfea8fe930042ff65ff11ff2c00370165ff30;
mem[606] = 144'h0147fdcd0108fe8a003b009d005f0009005f;
mem[607] = 144'hfeb0ff2bffbb008eff0bffe7feb4fde7fec5;
mem[608] = 144'hfac3fd6c018afcd7fecbfec70139ffa1004a;
mem[609] = 144'h014dff4effc6fffeff6d0109005302a30197;
mem[610] = 144'h043503ba03a702f3fe3f018904d305680412;
mem[611] = 144'hfe0200200120fc88ff97fc4a008efb79fc4e;
mem[612] = 144'h0109fc7f01ceff18ff1f00b20472001efe08;
mem[613] = 144'hffdeff2e013501d7fe4f012700fbff0a001f;
mem[614] = 144'hff4c003f0185fe2bfee800e1016dfea0fe37;
mem[615] = 144'hfdb6fea0fe28fe4efc4bfe4302e2026a01ce;
mem[616] = 144'h00ccfd3c00c70089ffb2004902b4023d0136;
mem[617] = 144'hff14fe8dfed4013b00d500cf01d401c6fe02;
mem[618] = 144'h01d8fb66012105eefd150002ff3ffb02fcad;
mem[619] = 144'h0086f85fffb10118feaa0084fb02facefd53;
mem[620] = 144'hfd66fcc8fe5dff3bfeb90434fe6afa20fda7;
mem[621] = 144'h037c04800344025cf929fb22078e0ea00d71;
mem[622] = 144'hfe2efebdfe0d0050010000fa00750050009c;
mem[623] = 144'hff1bff43fe86fff8ff27ffd7008e001eff7b;
mem[624] = 144'h0101fe16fe9200170143fddb006200bf0217;
mem[625] = 144'hffddfd67feae00b8014ffe9bfe28fdeafe86;
mem[626] = 144'hfe93002d012dfe5b00ebff3afdcb00a1016d;
mem[627] = 144'h0118feccfe3c01d7fee6fff7ff39fef90029;
mem[628] = 144'h01060080ff5e0103000a003401260081fe94;
mem[629] = 144'hff4dffc90022ff1fff6afec901b7ffbeff71;
mem[630] = 144'hfe89fe4fffc5fea5ffe6fde5fe940155ffc8;
mem[631] = 144'hff45ffe3ffe9fe4100d201270074008c0007;
mem[632] = 144'hfe9dff7500cc003b016f010fffa2015afdfd;
mem[633] = 144'hfe81fe64fe49ffedfe3000c9fd81ffa9fefe;
mem[634] = 144'h016fffa7015e006fffbb0249ffbdfe95ff55;
mem[635] = 144'h00bc0116fe53000a012200620034006a00e8;
mem[636] = 144'h0014ff300086005fffddfef40012ff08ffb7;
mem[637] = 144'hff2f0095ff2f002601b0ffef0128feaeff7b;
mem[638] = 144'h011cfe8bfec1fddd0120011ffea2fe19fe3f;
mem[639] = 144'h0038fe5d0112008dffd000190065ff4fffc5;
mem[640] = 144'hfd83fe0e00f90095ffcbffd1093600a1fe0c;
mem[641] = 144'h038dff19036bff6605300771048e02c802d4;
mem[642] = 144'h057604e9fddaff2a07380591008f06c40339;
mem[643] = 144'hfe1cfecbff9afd6affe6011c03a3ff15ff14;
mem[644] = 144'h0088ff65004802b5008e0128047f03b9fe6e;
mem[645] = 144'hfe660008fec8012600b8ffd2ff24fe4eff19;
mem[646] = 144'hfffdfe7a00b5009d0284053106dc02f0024d;
mem[647] = 144'hff40ff89fdeaff11fe1e0232035003410010;
mem[648] = 144'h0468fd8b0166ff30021a04da08e6060e0015;
mem[649] = 144'h067c00e5fef5feaa022e050e09ef054e00e2;
mem[650] = 144'h004cfdcefdb100c5fe5c0001fd0eff91fe12;
mem[651] = 144'hfd68fec3f8a503fefcfaffb1ff7f01abfb81;
mem[652] = 144'h0050ff42fe84f93bff7efdef022dfd60fe06;
mem[653] = 144'hfbc903050139031a009e022f00f5fdb800e0;
mem[654] = 144'h00c200f601f6fe81034e0626057e0225ff6f;
mem[655] = 144'h00e00028005cff17000c021c059f058f0184;
mem[656] = 144'hfe6cfebe003effff009c006bfeabff82012e;
mem[657] = 144'hffd6003eff0101c20096fe7800ba01f6feb9;
mem[658] = 144'hfeaf00a7fe37005600a1fe6fffa00185ffe2;
mem[659] = 144'hff6dff19fe05010cfe0bfdfcfdadff2bff4c;
mem[660] = 144'hfe550013fe86ffbdff210080ff1e0151fe49;
mem[661] = 144'hfe9a004ffef6fecc016500cb000dff6c01b1;
mem[662] = 144'hfe6fff1a012f00d2006b01160034003900b6;
mem[663] = 144'h007dffa100d3ff04fe42025700c5fec001c5;
mem[664] = 144'h003dffe5014b015fff150053ff9f00b7008b;
mem[665] = 144'h00f80096febdffeafffcff4801affd96ff4a;
mem[666] = 144'hffaffebcff6000ae0135ff63fe80fdddffba;
mem[667] = 144'hfef001310013001d00fdffdc00c7010ffe5d;
mem[668] = 144'hfda3fe0afffafe3efe86ff0f005d0156fe48;
mem[669] = 144'hfde0fe2d01a5005afdf1ffb2fec5febb0066;
mem[670] = 144'h01d6fe91ff0afdccff81ff5afeb7fe0d00e2;
mem[671] = 144'hffcf006c004c003efdd502540081fecc0080;
mem[672] = 144'h0138fe74fa6d01ac0435ff51012afb07fcad;
mem[673] = 144'h01d8fcf1f9e0037c0297011e01b8010c007a;
mem[674] = 144'h0059fc8506600752ff4500eb006407e1067f;
mem[675] = 144'h01f0ff66fc0605d703eefcc6fb40f992fb26;
mem[676] = 144'h02edfedcfc15fc6302c7032304ddff76fccb;
mem[677] = 144'h02120135ff8d0294fec7fe4ffe9fff80025e;
mem[678] = 144'h02cefe00fa02034a0609fef7fe86fae3fee4;
mem[679] = 144'h048802a6fd6afbd300a001aa0361fce4fcb9;
mem[680] = 144'hffb7fa97fde703150485032d01390191fff6;
mem[681] = 144'h039dfba5fbde002c05c4017e009bfce4fcf7;
mem[682] = 144'h01d004c109f2fa6eff6b026c023400eef9c2;
mem[683] = 144'h00ab04dd0262f954037a03ef0055fc48f4d1;
mem[684] = 144'hff54fd4dfb1508ec00c2fd5eff5afafefea9;
mem[685] = 144'h005207650608fdcf015f001802f208730159;
mem[686] = 144'h032ffb8df9e502f70657ff070020fe2a0192;
mem[687] = 144'h0346fe6bfcc9ffe10579027cfebffd69fd7d;
mem[688] = 144'hfddf0141035d0306fec4fd02006b02fc03ea;
mem[689] = 144'hffab038004200001fac901830089ffe8ff63;
mem[690] = 144'h00a700cc011afb85ff82022e0259fe45fc1c;
mem[691] = 144'hfde60183047802b1fc2b01a4004902220269;
mem[692] = 144'h01b001a000a10451fef2fed30132fedffe56;
mem[693] = 144'hfe11fdcfff28fd97fbbbfcf9fcddff68fd6a;
mem[694] = 144'h00f0ffdd059103defcdf0075fe8d005bff56;
mem[695] = 144'h014300b5014c059a0197fce5fed20193017a;
mem[696] = 144'hff5803cc0578ffcafe2cfe8f008bfd91fc42;
mem[697] = 144'h000d03dc048e035cfebdff440163ff9c00f9;
mem[698] = 144'h01f4feeef3eb040f04d2036d00df009bfe02;
mem[699] = 144'h031800b4fa57037b02f9fecb02c5019f01d6;
mem[700] = 144'h0230018f0467fc26fd290348004e0253037e;
mem[701] = 144'hff5cfce9fed9074e0272008fff3dfe5106ee;
mem[702] = 144'hfeae0114054b0101fecffffcffdf01530000;
mem[703] = 144'h00ffff5004220526ff8ffd2dffa50116019b;
mem[704] = 144'hff50053706b0062301b6fcd5004601acfff3;
mem[705] = 144'h026f031a016b017efd37fe9a0159fcbcfe19;
mem[706] = 144'h0090fa7bfb27fdb4fdb600b8fe26fc1cfec3;
mem[707] = 144'h03fa01c000170113fbbaff98027200a20111;
mem[708] = 144'h025c02300535016f0377fe930036ffdf0019;
mem[709] = 144'hfe020048fd8dfeddfd7bffb6fd68fef0fea1;
mem[710] = 144'h0392029503bd0088fd69007102f900d9fcb5;
mem[711] = 144'h0150ff32018502e102f201f2ff9101e60111;
mem[712] = 144'h00f003cc0014012b0169fec60221fdb40050;
mem[713] = 144'h00c603ca045b02870365fdbbffc0ff06fd39;
mem[714] = 144'hfe59f786f360fd0c01c3fed3fe79fdbffa25;
mem[715] = 144'hfd2efc06fc4dffb00352fe74fe00fe9dfc3b;
mem[716] = 144'h0285fe37fb64f891f89afee00205fb76fcf2;
mem[717] = 144'hff1efec4084303d40174fd3b0341035b049e;
mem[718] = 144'h030bffbbff2202b2fef8007c01e8ff0fff54;
mem[719] = 144'h0368032503c60284027201060057fe9c001a;
mem[720] = 144'hfb80fd8c00d5ff70fe39fcc9002a01b8ff2c;
mem[721] = 144'h0128011805e3fcf3fe0f02c4026002a2fd0b;
mem[722] = 144'h056808030068fc3a03bc03820390010ffc0e;
mem[723] = 144'hfac5fb360263fcddfee1005f02b6ffd10144;
mem[724] = 144'h00b8fc2cfce60209fe3efd1100a103ecfdb3;
mem[725] = 144'hfe41003e01f6011dfeef0193ff98ffd600ef;
mem[726] = 144'hfd57ff790263fe1afa7d00d1020b00f001b6;
mem[727] = 144'h00b4fdc3fdc50415ffc1fde3027404430193;
mem[728] = 144'hff460104025bfb04fdec005e04b70467fd4a;
mem[729] = 144'h0052fe96fe960013fb40fe92ffba0433ff82;
mem[730] = 144'h03b0001dfe8e097b0022016601ec054e0b71;
mem[731] = 144'hffb2feaefbb80638ff5ffd83ff3f04d9048f;
mem[732] = 144'hfff6febc05effbba02db02010454fead0349;
mem[733] = 144'h04fa01e5fb4404540112022e0076fe8a02d2;
mem[734] = 144'hfd2affbe01b9fe25fd50ffa7017f018e0109;
mem[735] = 144'hfd00fcc8ff8500dcfae9006002010403ff16;
mem[736] = 144'hff22feaf0098015500b8fe2d002e0122ffe9;
mem[737] = 144'hfffc009700fcff77feaafee3ffb300b101d5;
mem[738] = 144'hfde4fe36ffe7fe6c01dafe26fe4fff410169;
mem[739] = 144'h0028fee500010010fefc01c70044ff3b01cb;
mem[740] = 144'h006efec40015ffb20039ff4cffabfefffe55;
mem[741] = 144'h00590146fec10076fe59fe44feed001fff4f;
mem[742] = 144'h00a5ffc00002007c004bfebeff89ff0c00b2;
mem[743] = 144'hffea01b9010ffe93001cffbbfff500a300ee;
mem[744] = 144'h00e000ad011bfe5cff6700dc0032fe7cff1f;
mem[745] = 144'h0076fed3fe1aff27fdc5fff401bffe3cff83;
mem[746] = 144'h008bffe5ff3efe4efff7ffa200e6fedeff6c;
mem[747] = 144'h0002ff55ffafff06ff7b00cffe2d00a8ff87;
mem[748] = 144'h0056fff4015a01630029ff01ff1afedb006a;
mem[749] = 144'h00c7000f01defe9dff16ffcafed20099fe0d;
mem[750] = 144'hff0e00ca019f00a50013ff05ff2e00a7fe49;
mem[751] = 144'hfff5fe77fe37feebfe53007e013cfea80185;
mem[752] = 144'hfbeefd4b01ae018dfe0fffa40682037402da;
mem[753] = 144'h0337045a052a01ab03ab0681060f06110202;
mem[754] = 144'h062e09affff202bd072e048d046d0338fb9f;
mem[755] = 144'hfc31fe8302d1fcf5fbe7fd310574002504d5;
mem[756] = 144'h0392fe2cfecc0379ffb8ff8e0460046effde;
mem[757] = 144'h0163013a00b401a9016c0079ff40006c0051;
mem[758] = 144'hffa6003f05410080fecf03a605f7036b016b;
mem[759] = 144'hfe59fba5fea1032b004700fb034403750313;
mem[760] = 144'h0567026c053600d9041504ba06800571ffd3;
mem[761] = 144'h03a200d2033e0319021a04170748048e0208;
mem[762] = 144'hfff6fac5f61f04d4fc3100c5fd0bffe30270;
mem[763] = 144'hfdbff919f9780641ff1bff50ffef03b00190;
mem[764] = 144'hffcafed402f4f780fd54fd440292ff54001e;
mem[765] = 144'hfd66fe9bfd9c0276fecdff650210fe4f0784;
mem[766] = 144'h00a7fff306ba02be00430460038003f001e4;
mem[767] = 144'h0177006204a301d2ffdf010106a0036dffaa;
mem[768] = 144'h0144009afc9afddb00d60416008601c103ac;
mem[769] = 144'h0304010d048005c401690705fd73ff56ff4b;
mem[770] = 144'h01a6010906e6021d02e6021bff30fefbfa9b;
mem[771] = 144'h00280182fc83070702f7043e003c0224051f;
mem[772] = 144'hfde1013ffed4fd09ff1501d3fcf5fe63004e;
mem[773] = 144'hff26feab012dfeecfff900a0fea7fdc0ffdc;
mem[774] = 144'h0264007b029d03aa016304cf00af01b602cd;
mem[775] = 144'h0158020e00befea400ee032bfda400020268;
mem[776] = 144'h03c602d70232011501dc04befc9efdd60014;
mem[777] = 144'h0433035d01e002f100df03570025fe670203;
mem[778] = 144'h019507670b9efde2fda0fe82004208350553;
mem[779] = 144'hff8405ae0241fd9dff85019c0119084f05b3;
mem[780] = 144'h01bf05a1040604e2fd27ff7101f4048204d9;
mem[781] = 144'hfd20fd45f78bf5df030903f1ff4ffa3afb1e;
mem[782] = 144'h003900c801b4062c042005930070fe0effda;
mem[783] = 144'h0087037f021901e800fa04930176fffc03bd;
mem[784] = 144'hff3cfd7105dc0399ffc1fcc1010f013c0413;
mem[785] = 144'hff570195061afdadfca4003704a4020401f4;
mem[786] = 144'h03840453fc18fd2a0537026203f6012b015d;
mem[787] = 144'hfe94fdc704a2fe15fbce00530153017600dc;
mem[788] = 144'h009400ca017906b5007afeaa044b00e6017d;
mem[789] = 144'hfe9e008eff35fff7ff110140fe5bfd78fd43;
mem[790] = 144'hffd0ff5e049e015dfb3efee8021c02270181;
mem[791] = 144'h00c6fc5f018803d0ff01fdb5037c01100058;
mem[792] = 144'h004a015204a300ab000100a5048cffc5ff9b;
mem[793] = 144'h000300a5050b0365fde0fec3038b032e01eb;
mem[794] = 144'hff42fb21f47704f305a00043fdd6fdf6fb74;
mem[795] = 144'h0330fb0ff835052002f3fd200149fee2fcdc;
mem[796] = 144'h0101ff0a0291f6e8fbf503c10423001c0151;
mem[797] = 144'h0052fe76057e0ba8fd6fff0400fb02ce05ef;
mem[798] = 144'h01da0134042a01d2fbb0fe81036d00520361;
mem[799] = 144'h003100d803b702310008ff9b028b011b0205;
mem[800] = 144'hfde0ffdb0171fe710030fea9ff3a00490043;
mem[801] = 144'hfef3ffa4009c00f8fec100a7002eff1e011d;
mem[802] = 144'hff95fe65fe22ff7afeec0055feb1ffa600ad;
mem[803] = 144'hfe29016c0067fd20fecb01580072fe55feec;
mem[804] = 144'hfe0affeeff80006ffe4eff1c007000e4fd97;
mem[805] = 144'h0057ffe0fe3b0017ff02ff96ffcc006d0121;
mem[806] = 144'h008900b9ff58ff7c008100e0ff910189fef9;
mem[807] = 144'hff94ff6e0023006900f0fe0afe4fff22007f;
mem[808] = 144'h00c900be004aff32fe7afdbbff1cfee200e1;
mem[809] = 144'hfeac0080fecafefcff47fe72fea2ffb400c8;
mem[810] = 144'h0090007dfda30058fd2efd4ffe51fdb8ff97;
mem[811] = 144'hfec0fec2fea9009bfd6efdc9fe32ffeffd2d;
mem[812] = 144'hffd2fda4ffddffde00bfff27fea6feef0003;
mem[813] = 144'hfff100e2ff47fe03fe5efec5ffb7019ffe39;
mem[814] = 144'hff43fe07fdfbfed0ff4cfe7efe8bfe8eff99;
mem[815] = 144'hfe81ff3ffefffe47ff040033fd61fe94ffad;
mem[816] = 144'hffa4fdd4fbbaff78036801d5ff8dfb7bfee2;
mem[817] = 144'h00cafb7cfd7b021c031400c60161004804db;
mem[818] = 144'h008a02ff05fc001afe41006802570561036d;
mem[819] = 144'hfd0bfd2cff320407043100eafdd0fe320042;
mem[820] = 144'h0075fd9efb31fe250366055f019500b3fc65;
mem[821] = 144'h00edfebeff1702df01a6ff970143ffedfefa;
mem[822] = 144'hff6ffbf1fe4b00b40164fec901ddfe95ffbd;
mem[823] = 144'h01c700e0fa21ffa3011502a30433fd85fcf0;
mem[824] = 144'hfcf0fd3efd4b00ef0156000701d3ff4f0134;
mem[825] = 144'hfd34fc22fc12ffbe0134024b03f6ffeefe6f;
mem[826] = 144'h02a109f105b2fd41fd3c01fcffc401b4f9bf;
mem[827] = 144'h037007affa00ffddfeaa0373004000d4f86a;
mem[828] = 144'h013afda8024304980480ffeeffd0fe4e0184;
mem[829] = 144'h023d0483ff2d000f0069012f036f046100cb;
mem[830] = 144'hff0afbd3fc0a01430396fde6ff5eff83023c;
mem[831] = 144'hfe2afc7ffb38ff3403710310001a002c00d2;
mem[832] = 144'h000e01c000c6025000c1025bfa1e00c303f2;
mem[833] = 144'hfa9d03a30375fcedfbbefbbdfb78fd5eff87;
mem[834] = 144'hf930fe900275f9d8fb59fa28ffaff35cfb22;
mem[835] = 144'h044405040140ffff024302e5ff6a050002df;
mem[836] = 144'hfcfa0210039d014ffdf7fe9df7ebfc72012e;
mem[837] = 144'h01c203f800a1003c020700edfe6cffe10089;
mem[838] = 144'hfea602f602b60065ffa2fd9ffc030123fe45;
mem[839] = 144'hfe58023504ee00d9fea00008fb9d01b8ff47;
mem[840] = 144'hfa3204930497ff53fd2ffcc7f983fe85018d;
mem[841] = 144'hfc08044e010dfd27fe5efdd0f877fde5ff14;
mem[842] = 144'h023803be0478ffdf04d5038105f00125094b;
mem[843] = 144'h02540509053801e500b50351031700e7092d;
mem[844] = 144'h01e108ba00af001003600105fe9d066d0321;
mem[845] = 144'h039ef719f95901b104c1015efe08ffb5febf;
mem[846] = 144'hffab032c004dfeb0007efd55fc1dfe48fd27;
mem[847] = 144'hff72017d000700cd00cafed4fcbc011b01e5;
mem[848] = 144'hfdbcfd53fb59fd4b00700547010c016d0231;
mem[849] = 144'hffddfd53fd66027402ed00f2017f046903fb;
mem[850] = 144'h020a03c105d40920019601190066032504a0;
mem[851] = 144'hfdd3fe3efc1400a602f00100014fff570339;
mem[852] = 144'hfed3fc4afae1fc83007304e5fe2b02c2030f;
mem[853] = 144'h01e9022100b9028f0375022d0309024e01fb;
mem[854] = 144'hfd7dfd6bfe03015603ff045dfeb10242062d;
mem[855] = 144'hff06ff6dfecbfd93fd8f0497000000410457;
mem[856] = 144'hff67fc33ff01021804240311fd220507043c;
mem[857] = 144'h0045fdd6fb0f001e01e9042c00c601fb0325;
mem[858] = 144'hffd10a1b122afffbfbd8ff88fe98ff48f9d0;
mem[859] = 144'hff6502ad0421fdf5fd83020e002ffea80284;
mem[860] = 144'h015500b9035206b2051c0104ffa600ad00d7;
mem[861] = 144'h031f022ffb98f3bbfc2dffc1038bfed3fc51;
mem[862] = 144'hfdc4fedfff1901a205760118ffa3021e036b;
mem[863] = 144'hfe28fc5ffde5ff8a01c7024afe9c02f1040d;
mem[864] = 144'h02f9024ffd69fcc6ff1904e80448ff52ffdc;
mem[865] = 144'h04ba0135f8a1ff8e014501fdffbf02070475;
mem[866] = 144'h024efcf8fe53057f00a1ff62fc920007053e;
mem[867] = 144'h03b400f8fbcbff58038804e0045400500101;
mem[868] = 144'h00e400a802b9fa7efbfb033e013102940212;
mem[869] = 144'h0273ff2b016402f900bb018902d603d4040a;
mem[870] = 144'h012c02ddfc4dfff7036606950319021f012d;
mem[871] = 144'hfd9304900244f958ff1b01780119020f00f3;
mem[872] = 144'h03030110fda201c9006b02e3004f020f0554;
mem[873] = 144'h02cb0184fee7ffb6ffbc045d0138031e0615;
mem[874] = 144'hff0903cb0be70388fe97fba5fe7003cbfe73;
mem[875] = 144'hff450093068efe42fb1bff8e0025041901ee;
mem[876] = 144'h041e005d005e061701c50028010f03b801cc;
mem[877] = 144'hfb9ffde8fd26f5c8fb5402adfee7fc4af60a;
mem[878] = 144'h023d028ffc6efd67038c0669048101e8037a;
mem[879] = 144'h03c701d0fe32fe50001803cd04b500fe0303;
mem[880] = 144'h00c300f4fd72fd71fef2ffbc0489ff0c0309;
mem[881] = 144'h029afec3fcfb025e0117ffd1039204520550;
mem[882] = 144'h00300022008c0396fe8e008cfe120679020c;
mem[883] = 144'hfe72fde0fc1602640115fe3001fbffc3011a;
mem[884] = 144'h0018ff3c01feff4d001bfe4a03ab02b701bb;
mem[885] = 144'hff83fd4b00acffdefffbff0301a2fdfffd3d;
mem[886] = 144'h04370119fef900e602f401d904130100028a;
mem[887] = 144'hfea5003bffc1fe9a00d4007d00ed021f0004;
mem[888] = 144'h05740011fe270068fef5ff3204e3052b0254;
mem[889] = 144'h03d500bbffd2fff2ff1101e7051402310483;
mem[890] = 144'hfff1fdc5fdc6011afe38fefaff43fd38f7f3;
mem[891] = 144'hfffdfa52fc40fd0dfdc4ffb9ff280166ff49;
mem[892] = 144'hfecbfd6f009d0173fcacfc9cff880135004a;
mem[893] = 144'hf8c30299fe6ff93efd92007dfedef96afc81;
mem[894] = 144'h0302ff81006e013803ad034c040603630493;
mem[895] = 144'h02110138fec4017a01c5ff3a061c006b0523;
mem[896] = 144'hfe09fb50fddfff64fb4cf86bfc5301aa01e5;
mem[897] = 144'hfe9100c8039fffe9fce5fac500aa002d01c6;
mem[898] = 144'h0395050708a7022dfeee0249030002820030;
mem[899] = 144'hfe48ff8c002a01bffcedfb5b0003005c002c;
mem[900] = 144'h00630018fbc8ff14fe23f93dfde900cdff88;
mem[901] = 144'h00e401f302750219007300c3011a00d80151;
mem[902] = 144'hfe05fc6201d8ff37fb31f72bfd1302210075;
mem[903] = 144'h0165fdabfe0cfff6fe4df99dff7f016a0053;
mem[904] = 144'hfe7d026c0324fe54f9c7f9edfe3002a80038;
mem[905] = 144'hfdbbfe06ffc2fe51fd28f951fc0a0250feb2;
mem[906] = 144'h048806b304aa069d040000e701bffcdc0595;
mem[907] = 144'h031401f3fe6f02ec001afedaff5afef102ee;
mem[908] = 144'hfebf0262028202d4011c069900a40165ffc9;
mem[909] = 144'h02e50187fb9cfecdfed5ff940389067902b2;
mem[910] = 144'hfd97fde90175ff21fe69f7dcfdc002bcff1c;
mem[911] = 144'hfcefff79fda4fe0cfdb6fa5ffe64028600c4;
mem[912] = 144'h011ffe29ff74fe4400ebffbdff05ffab010c;
mem[913] = 144'hff37ff370006fe2cff6bfe7dfe70ff680057;
mem[914] = 144'hff77fd7d00bbfd9c00f100a600ddfec00123;
mem[915] = 144'h00000047000b000900c3fe70ff42fe7bfde8;
mem[916] = 144'hff5e0007ffcbfff9ffc8fd9dfda900f1fe4d;
mem[917] = 144'h006c01d2fe5bfe7600a7ff4cff59ffe50126;
mem[918] = 144'hfeab009dfd7e0074ff320029fee3ff5efdfd;
mem[919] = 144'hfec7fdbcffe5ff360027011cffd5fd9b00d9;
mem[920] = 144'h00900050fe23ff65fe00fe1200c1fefafdf9;
mem[921] = 144'h000f0078ffdcfe7afe5cfeebffeefee5fd70;
mem[922] = 144'hfe1eff09fdfdff78ff470116ff77ff49ff24;
mem[923] = 144'hffe6fffdfe61fe1ffed3002e01c3006dfdc0;
mem[924] = 144'hfd82ffd70199fe96feeefff7ff8dff8dfd88;
mem[925] = 144'hff4bfefc0065fe0cff54fefffda9009f0087;
mem[926] = 144'hfeaefe26fdf1fde3ff8a00a7fdcaff78fffc;
mem[927] = 144'h008f006b008efda6fe72ff9d003c0016ff3b;
mem[928] = 144'h015a050e02d8026c01c700dafbf9036e029b;
mem[929] = 144'hfe5805f504430325fb11fc49fcefff16fba8;
mem[930] = 144'h003001bcfe41f88cff31ff82fe79f4c2f762;
mem[931] = 144'hffc90161ff05030cfba3ffe201af05150152;
mem[932] = 144'hfeb004c2014aff6f033bfdacfc2ffd21004f;
mem[933] = 144'hfebbff0dffd8fcdbfde10033fe5dffe8fe7a;
mem[934] = 144'h00c601a001580338ff2cfbb4fc0100e50161;
mem[935] = 144'hfea8030d021d00dd0130fed5fc6aff27ff4a;
mem[936] = 144'hff1204b900790024fe95fdbdfa1afcca0052;
mem[937] = 144'hfef0041a0159031c016dfd0bfc56fd21fff5;
mem[938] = 144'hfff7fb19fb55f97f028800a80279041d07cc;
mem[939] = 144'hfe79fe31018afd9704ad01ee003203df0645;
mem[940] = 144'h016a041101e0fca5fb03fffe003a0430fe87;
mem[941] = 144'hff46fb6ffd0200d9074305abfcadfccffc2f;
mem[942] = 144'hffc404500261ffbdfcd0fc34fe7bffd7fe6c;
mem[943] = 144'hff40031b02aa02e6ff70fc0cfbff000dff5c;
mem[944] = 144'hff50003b00fcfdb90121fd7dff960047fd87;
mem[945] = 144'hfe1c0031ffc3fdc6ffce00f0ffc4ff15ff69;
mem[946] = 144'hfed8febc0024fe86002a0062ff26ff6cfe1e;
mem[947] = 144'hfd8c005ffe9d004dfd9bfe89ff0b0096fdd8;
mem[948] = 144'hffefff6c002efe64ff31000dff03ffa2ff8d;
mem[949] = 144'h008f006f014400d001aeffe100d0fe8fff92;
mem[950] = 144'hfefcfffb00eaffe600820106fe310075fdd1;
mem[951] = 144'h000a00870000fdd8fdc3fe740051ff7dfeeb;
mem[952] = 144'h00f4ff4bffc2ff10ff53ffb8fe360061feb7;
mem[953] = 144'hfe73ffc2fe25fdceffe8fd9aff1affcafe49;
mem[954] = 144'hff0e0096fd8ffd95ff83ffd300310118fd99;
mem[955] = 144'h002a0000fe420092ff240070feaf0073ff75;
mem[956] = 144'hffbffe23fe59fdaafe830025fd90fff000b8;
mem[957] = 144'hfe59ffdcfe00ffe1fdc4fe27ff94fdadfe2f;
mem[958] = 144'h003500e4fe23fe5a00c1fe88fe07004ffe33;
mem[959] = 144'hff7a00a7ffecfff6ff3ffe96fe1500defdbc;
mem[960] = 144'hfde4012dfea9fec8ff5e0163ffedfff4fe4e;
mem[961] = 144'h01d700200043fed0ff25feb6fe2fff5affb7;
mem[962] = 144'hfebefeac017201bf00e100cf001100400023;
mem[963] = 144'hff62ff3d0066fe46fe98ff55fee10154feed;
mem[964] = 144'hfe59fe71ff56ffa8fe42015b0144feb3fefe;
mem[965] = 144'hfef600b7fec301b80053febb0129fecbfef4;
mem[966] = 144'h002d011fff18fdef00c1feb0fffc002d00f9;
mem[967] = 144'h0163ff8f01050127fe89fe9cfeabfe64ff21;
mem[968] = 144'h0018fee3fe3dfe6eff7fffdd0055ffe00118;
mem[969] = 144'h0180fffa0144ff8e000f006200a000a4017e;
mem[970] = 144'hfe97fdda0165010dfe9f0155fe5bfdf5ff01;
mem[971] = 144'hff86fe09ff63ff02004eff12001d0137ffdd;
mem[972] = 144'hfe01fe86ff52009d0035007effffff8cfe62;
mem[973] = 144'hfe2800c0fe13ff09fec5fff2ff5e00a5fe62;
mem[974] = 144'hfebdfde4ff1d004cff23fe2ffe24fecc004a;
mem[975] = 144'h015fffe3ff5000b2fe47fe200035ffb9010b;
mem[976] = 144'hfd4dff73ff09fde1fdfffff9fd24ff01fde0;
mem[977] = 144'hfd37022e031c025b0061fd96ffe1fd40fd8f;
mem[978] = 144'hfe15008d0046003d0080ffabfffffd65001b;
mem[979] = 144'hfd2fff6ffe7d0298ff9300adfcb80019ff43;
mem[980] = 144'hfffdfd12001efe77ff39fe9ffdd9fcd6ff2b;
mem[981] = 144'hff9d001800adfe970023018e0124ffaaff19;
mem[982] = 144'h00290268fe5ffdc10045fd7d0017fe3afe85;
mem[983] = 144'hff7300b90097fe260063003900c40148fda4;
mem[984] = 144'hfe9bffbb0257fd01fceb006afe3fff0bfef1;
mem[985] = 144'hff03030e00befe29fd1cff89001dfd14ffbd;
mem[986] = 144'hfef00001ffd400b80030001ffe44007b004a;
mem[987] = 144'hff77ffd80012ff48ff2ffcf3ffd6fe2ffdbb;
mem[988] = 144'hfe11fe9cfda700620071fe5bfd59fd7bfd22;
mem[989] = 144'hfd49fdcfff23fd51fe14fd6efed0ffe400b5;
mem[990] = 144'hfe9fffae031a00b1fd2c0078fd1ffd5efce6;
mem[991] = 144'hff700241005b0073fd16fe71fcd9fe85fdfa;
mem[992] = 144'h02d901e403d4050dfef2fe44007cfe3700e2;
mem[993] = 144'h025c002c0066036d02300340ff56fe8c0026;
mem[994] = 144'h01a9fddcfaf5fed704ba02460004027efc63;
mem[995] = 144'h001cff7e037d0029fc1e03c3ffd5fd570487;
mem[996] = 144'h0491ffb8ffb004a802a50104026dfe74fef4;
mem[997] = 144'hfd02ffcffd340025fe60010200a5fc9ffd5f;
mem[998] = 144'h042f0191015203f2fdf0030d0110ff37019b;
mem[999] = 144'h047302d0ff6c0343010801d602dffeea0027;
mem[1000] = 144'h040a0120026b0407032101f3023e00e1fe0a;
mem[1001] = 144'h0397ff30027d0556006603e7042f0047feaa;
mem[1002] = 144'hfe52000af4a70289ff870057ff2002cff9b5;
mem[1003] = 144'h0062ff31f8ad03d9ff0eff9affe20271facf;
mem[1004] = 144'h0322fe1105abf99cfcc5ffe3ffcdff51046d;
mem[1005] = 144'hfe9100b10122008b017cfe9403acfe390170;
mem[1006] = 144'h0336009701330407fe3d032affea013e01f2;
mem[1007] = 144'h04bc00c903a2059100340355043001610269;
mem[1008] = 144'h016300dffd61ffc101c2ffeefd13fc78fbe6;
mem[1009] = 144'h000cfce2fea90098ffbefe360139ff380116;
mem[1010] = 144'h0079fe85091104fefd73012e01ff08b9071d;
mem[1011] = 144'hfd30fd9dfcd70320026dfbcffb9efc05fe72;
mem[1012] = 144'h013dfecffed6fe030206009f009b000fff42;
mem[1013] = 144'h0055002203730055fe0fff0cfe81024d0178;
mem[1014] = 144'hfe0bffd5fed3feb503a9fdbcff18fc6e0078;
mem[1015] = 144'hffa3febbfeb8008d001e018f010ffeb8ff92;
mem[1016] = 144'hfbc8fdf1fc9afed4fe6600b2ff76fe9a0132;
mem[1017] = 144'hffcdfe1afd5600b8023dff160053ff9efd6e;
mem[1018] = 144'h0328018900c501150363001f015dfb90fa67;
mem[1019] = 144'h01f0fe3701fbfee30189009c00edf998f99f;
mem[1020] = 144'hff51fbf3f9e508070146049bff85fcf00123;
mem[1021] = 144'h010e025702b0ffd80027feea0276050a038c;
mem[1022] = 144'hffdcfd8afcbe025801cffe89ffa3fda2ffc8;
mem[1023] = 144'hfdf2fd6dfc8cfec40264ff26ff3afc7dfe45;
end

always @ (posedge clk) begin
	q_a <= mem[addr_a];
end

always @ (posedge clk) begin
	q_b <= mem[addr_b];
end

endmodule