`timescale 1ns/1ns

module wt_mem2 #(parameter ADDR_WIDTH = 11, DATA_WIDTH = 144, DEPTH = 76) (
input wire clk,
input wire [ADDR_WIDTH-1:0] addr_a, 
input wire [ADDR_WIDTH-1:0] addr_b, 
output reg [DATA_WIDTH-1:0] q_a,
output reg [DATA_WIDTH-1:0] q_b
);

reg [DATA_WIDTH-1:0] mem [0:DEPTH-1];

initial begin
mem[0] = 144'h05bfe1c3fa4607781b81fc08086cf6b50ecf;
mem[1] = 144'h0584297f0b7327d50f6008281b7d0177fdfd;
mem[2] = 144'h012e00ec006308b8059e0cb1fd71f9d608ae;
mem[3] = 144'hf72b001a026dfe170ae008a3f86c00d2042a;
mem[4] = 144'h06510437fe8f0314084407d8ff4af7a0fdc3;
mem[5] = 144'hf6b5fc1a091cfaf2058304caf81601a701f3;
mem[6] = 144'h068afe2f00cf036d04ab07adf9bcfbad0d27;
mem[7] = 144'hfda903d9042804490e8e00f5f8c5020103b6;
mem[8] = 144'h0b700a53fa870aabffeafa2c08000420fe3f;
mem[9] = 144'hf801f0c6f663fbdaf56400f703ef056f0966;
mem[10] = 144'hfe60ef52f43ee8c3de14e92bf425f391f0bc;
mem[11] = 144'hf202eb56fbedee83f0fc043cfb1d049e0fdd;
mem[12] = 144'hef07f9fdf3880504fd3100c705220d980c19;
mem[13] = 144'hfe06f54df609fd22fc55fe36007100c30a5b;
mem[14] = 144'h01b6020ef56505fbfc140152ff19fb1dfb31;
mem[15] = 144'hf793f6120397fb210aab0ca2077c0451fc52;
mem[16] = 144'hef95e6a9f28cea9adba8f4dcede1f434faf1;
mem[17] = 144'hf81ef51e08f0ed0efdbb106afd750adb005f;
mem[18] = 144'h08c6053dfce40356fc0f04e7fc86f84c007e;
mem[19] = 144'hfa5efe680418f707038e05f5015c05d207a5;
mem[20] = 144'h05df01ec020b074808e80ce4fb4705c810ce;
mem[21] = 144'hfbbafe1dfae0086a0c67fb64fd3fff7bfa96;
mem[22] = 144'hf156f41beed1ef79f14feac5f4920068f1de;
mem[23] = 144'h074206e8002412030816f956108e0a99f39e;
mem[24] = 144'hfb200145fe85013cfad402bfffb5fcc2fdbf;
mem[25] = 144'hfcbdfa87fd8dfaf8fd56fce4fe34fdc502df;
mem[26] = 144'h039b046bff6c16fc0a1efe5f12eb061efb57;
mem[27] = 144'hfb12f022ee61f893fcc2f6eeff54fe380540;
mem[28] = 144'hfa500476f8c9f744f0f6f250f8edfbccffc2;
mem[29] = 144'hf15a0062060efa3e07ac09ed026806a3fd82;
mem[30] = 144'hf902f5eff198f6b2f0b1f3e5ff93097efdf4;
mem[31] = 144'hfc9eedabf6baf885f624fc31ffda002705d8;
mem[32] = 144'hfdbbfd5bfa03fcd0088f09e6f35c006609e7;
mem[33] = 144'hfda6fcd60260fecf040801d0fff105e1fa26;
mem[34] = 144'h0a2c07ba00a5028d057b04ccfbd500970bc7;
mem[35] = 144'hf306fe5af9ddf7e807d30cf6f735fbea0150;
mem[36] = 144'h0622012d01270a2a04c9fa8c0b74055b01a8;
mem[37] = 144'h02c2fcd5faa0ffc3f92d0119fffafe600919;
mem[38] = 144'h0b4812ea07180f8616c117ccfb8b079a0b33;
mem[39] = 144'hf8acfa0cf4c401a5093e06fef2c20912fc82;
mem[40] = 144'h0e020b2407910c7507a501c8fad9f9e804f3;
mem[41] = 144'hf410fc3201dafce502d80210ffa811d80b20;
mem[42] = 144'h03cb016afc7401fa008204e4f8d3fa8a030f;
mem[43] = 144'hf83efbfffc1102fe081d017dfcd109ef0489;
mem[44] = 144'he6a8ec42f825ea3df645f231f320f9f9f7d7;
mem[45] = 144'h09eb0725fa6c0839040ff61605bb0071eed1;
mem[46] = 144'hfc33e147e9c0f56fe11ded28ec84dbb3f0b0;
mem[47] = 144'hfd19f4910321f88df35e0ac9ecd9f9f50971;
mem[48] = 144'hed61ec45f22ff81cfcecf752f4a403cf02ea;
mem[49] = 144'h0aa30eb8fce108420aa0f28c03660a81f689;
mem[50] = 144'hfc3b03e7043c00d6fc4ffc08fd85feebfc8c;
mem[51] = 144'h0078ffc300f4002d02e703a00286f9f8fe99;
mem[52] = 144'hf5a2e744efcbfbcae17ae1f5e9b8d6a0ed94;
mem[53] = 144'hff60f405fc50f9d5f1a30420ee88fd410d73;
mem[54] = 144'hfd8f0536020804e201f0fdd80530012501e4;
mem[55] = 144'h02fc03a603e9fbb500e5fd15022bff7604fd;
mem[56] = 144'h123f0f7417d60173016b0679019df8c6f6d7;
mem[57] = 144'h0f220c180d37044809760291f412ef3de8bb;
mem[58] = 144'h00e7031e087108bf103211f6f845ffc20acf;
mem[59] = 144'hfa170d69051506f107c80bb6f4daf943f815;
mem[60] = 144'hf880ff75fa7bfecbf9eaf884fbf3fbcef9f0;
mem[61] = 144'hf085fb17fbd8f94a02b601a8fed004280010;
mem[62] = 144'h01c40479fa21050b04450672f59301a406f5;
mem[63] = 144'hfb3f02ed0266046f0b9d0471fabd055901a6;
mem[64] = 144'hfedd0010f4b2006ff9f7fa20fc7ef6d106ea;
mem[65] = 144'hf81202cf0491f958093c034ffc61066f0230;
mem[66] = 144'hfd1cf9f00398f88804d40392f6f0fb990046;
mem[67] = 144'h00f500420301fdda05b7fd2302b40345f83b;
mem[68] = 144'hfae3fdd6f7d1f875094306e10654077afde9;
mem[69] = 144'h04a30602ffbbff14ff5e05c9ff93fea30224;
mem[70] = 144'h0661f9a4089f0af306d6fa17f92509d0ffe6;
mem[71] = 144'h0737fc27f94102eb0428f9baff4606fe0233;
mem[72] = 144'hf892fa71023f0545fda7fad8fa85f59bfaef;
mem[73] = 144'hf96b0470fd3a0314fd9402a5fcf007fefeea;
mem[74] = 144'h0673f87af6b50528f76f0221fc47f1b7f8f8;
mem[75] = 144'h03e7fe41023cfd36fc1f02db056e07b9024d;
end

always @ (posedge clk) begin
	q_a <= mem[addr_a];
end

always @ (posedge clk) begin
	q_b <= mem[addr_b];
end

endmodule