module CNN_test
(
    input clk,
    input rst,
    output [7:0] pixel_i,
    output pixel_i_valid
);
    logic [30:0] count_time;
    logic [3:0] digit_w, digit_r; //state
    logic [4:0] x, y;
    


    //counter
    Counter #(
        .WIDTH(30),
        .MAX_COUNT(50000000)
    ) counter (
        .clk(clk),
        .rst_n(rst),
        .enable(1'b1),
        .count(count_time)
    );

    //digit
    Counter #(
        .WIDTH(4),
        .MAX_COUNT(9)
    ) digit_counter (
        .clk(clk),
        .rst_n(rst),
        .enable(count_time == 30'd49999999),
        .count(digit)
    );

    //xy  
    Counter #(
        .WIDTH(5),
        .MAX_COUNT(29)
    ) x_counter (
        .clk(clk),
        .rst_n(count_time == 30'd49999999),
        .enable(1'b1),
        .count(x)
    );
    Counter #(
        .WIDTH(5),
        .MAX_COUNT(29)
    ) y_counter (
        .clk(clk),
        .rst_n(count_time == 30'd49999999),
        .enable(x == 29),
        .count(y)
    );

    //pixel

    logic [29:0][29:0] digit_1 = '{
            30'b000000000000000000000000000000,
            30'b000000000000000000000000000000,
            30'b000000000000000000000000000000,
            30'b000000000000000000000000000000,
            30'b000000000000011000000000000000,
            30'b000000011111111000000000000000,
            30'b000000000000011000000000000000,
            30'b000000000000011000000000000000,
            30'b000000000000011000000000000000,
            30'b000000000000011000000000000000,
            30'b000000000000011000000000000000,
            30'b000000000000011000000000000000,
            30'b000000000000011000000000000000,
            30'b000000000000011000000000000000,
            30'b000000000000011000000000000000,
            30'b000000000000011000000000000000,
            30'b000000000000011000000000000000,
            30'b000000000000011000000000000000,
            30'b000000000000011000000000000000,
            30'b000000000000011000000000000000,
            30'b000000000000011000000000000000,
            30'b000000000000011000000000000000,
            30'b000000111111111111111110000000,
            30'b000000000000000000000000000000,
            30'b000000000000000000000000000000,
            30'b000000000000000000000000000000,
            30'b000000000000000000000000000000,
            30'b000000000000000000000000000000,
            30'b000000000000000000000000000000,
            30'b000000000000000000000000000000
    };

    logic [29:0][29:0] digit_2 = '{
            30'b000000000000000000000000000000,
            30'b000000000000000000000000000000,
            30'b000000000000000000000000000000,
            30'b000000000000000000000000000000,
            30'b000000000111111111111000000000,
            30'b000001111000000000000110000000,
            30'b000110000000000000000110000000,
            30'b000000000000000000000110000000,
            30'b000000000000000000001100000000,
            30'b000000000000000000111000000000,
            30'b000000000000000011100000000000,
            30'b000000000000001110000000000000,
            30'b000000000000011000000000000000,
            30'b000000000000110000000000000000,
            30'b000000000001100000000000000000,
            30'b000000000111000000000000000000,
            30'b000000001110000000000000000000,
            30'b000000001100000000000000000000,
            30'b000000011000000000000000000000,
            30'b000000110000000000000000000000,
            30'b000001100000000000000000000000,
            30'b000001100000000000000000000000,
            30'b000011111111111111111110000000,
            30'b000000000000000000000000000000,
            30'b000000000000000000000000000000,
            30'b000000000000000000000000000000,
            30'b000000000000000000000000000000,
            30'b000000000000000000000000000000,
            30'b000000000000000000000000000000,
            30'b000000000000000000000000000000
    };

    logic [29:0][29:0] digit_8 = '{
            30'b000000000000000000000000000000,
            30'b000000000000000000000000000000,
            30'b000000000011111111100000000000,
            30'b000000001111111111111100000000,
            30'b000000111111111111111110000000,
            30'b000011111000000000001111000000,
            30'b000111100000000000000111110000,
            30'b000111100000000000001111100000,
            30'b000111110000000000011111000000,
            30'b000001111100000000111100000000,
            30'b000000011110000011111000000000,
            30'b000000000111111111100000000000,
            30'b000000000011111110000000000000,
            30'b000000000111111111110000000000,
            30'b000000000111100011111000000000,
            30'b000000001111000000011111000000,
            30'b000000111110000000000111100000,
            30'b000001111000000000000001111000,
            30'b000011110000000000000001111000,
            30'b001111000000000000000011110000,
            30'b001111000000000000000011110000,
            30'b000111100000000000000111100000,
            30'b000011111111111111111111000000,
            30'b000000111111111111111100000000,
            30'b000000001111111111100000000000,
            30'b000000000000000000000000000000,
            30'b000000000000000000000000000000,
            30'b000000000000000000000000000000,
            30'b000000000000000000000000000000,
            30'b000000000000000000000000000000
    };

    assign pixel_i_valid = count_time < 30'd901 ? 1 : 0;

    always_comb begin
        digit_r = digit_w;
        if (count_time == 30'd1000) begin
            case (digit_r) 
                4'd0: digit_w = 4'd1;
                4'd1: digit_w = 4'd2;
                4'd2: digit_w = 4'd8;
                4'd8: digit_w = 4'd1;
                default: digit_w = 4'd1;
            endcase
        end
        case (digit_r)
            4'd0: pixel_i = digit_1[y][x] ? 8'hff : 8'h00;
            4'd1: pixel_i = digit_2[y][x] ? 8'hff : 8'h00;
            4'd2: pixel_i = digit_8[y][x] ? 8'hff : 8'h00;
            4'd8: pixel_i = digit_1[y][x] ? 8'hff : 8'h00;
            default: pixel_i = 8'h00;
        endcase
    end

    always_ff @(posedge clk) begin
        if (rst) begin
            digit_r <= 0;
        end
        else begin
            digit_r <= digit_w;
        end
    end


endmodule