// node structure: https://www.researchgate.net/publication/317574806_Automated_Systolic_Array_Architecture_Synthesis_for_High_Throughput_CNN_Inference_on_FPGAs  

