module num2pixel(
    input[3:0] num,//0~9 : 0~9, 10 : =, 11,12,13,14 : +-*/
    input[7:0] addr,//'d0~'d99
    output[9:0] brightness
);
    logic [7:0] asciipixel;
    assign brightness   =   {asciipixel,2'b00};
		if (num == 'd0) begin // 0
			case(addr)
				8'd00:asciipixel = 8'hff;
				8'd01:asciipixel = 8'hff;
				8'd02:asciipixel = 8'hff;
				8'd03:asciipixel = 8'hff;
				8'd04:asciipixel = 8'hff;
				8'd05:asciipixel = 8'hff;
				8'd06:asciipixel = 8'hff;
				8'd07:asciipixel = 8'hff;
				8'd08:asciipixel = 8'hff;
				8'd09:asciipixel = 8'hff;
				8'd10:asciipixel = 8'hff;
				8'd11:asciipixel = 8'hff;
				8'd12:asciipixel = 8'haa;
				8'd13:asciipixel = 8'h2b;
				8'd14:asciipixel = 8'h3;
				8'd15:asciipixel = 8'h0;
				8'd16:asciipixel = 8'h7;
				8'd17:asciipixel = 8'h3c;
				8'd18:asciipixel = 8'hc9;
				8'd19:asciipixel = 8'hff;
				8'd20:asciipixel = 8'hff;
				8'd21:asciipixel = 8'hce;
				8'd22:asciipixel = 8'h4;
				8'd23:asciipixel = 8'h85;
				8'd24:asciipixel = 8'hc8;
				8'd25:asciipixel = 8'hcc;
				8'd26:asciipixel = 8'ha2;
				8'd27:asciipixel = 8'h1;
				8'd28:asciipixel = 8'h13;
				8'd29:asciipixel = 8'hf1;
				8'd30:asciipixel = 8'hff;
				8'd31:asciipixel = 8'h7d;
				8'd32:asciipixel = 8'h47;
				8'd33:asciipixel = 8'hff;
				8'd34:asciipixel = 8'hff;
				8'd35:asciipixel = 8'he2;
				8'd36:asciipixel = 8'h20;
				8'd37:asciipixel = 8'h30;
				8'd38:asciipixel = 8'h16;
				8'd39:asciipixel = 8'haf;
				8'd40:asciipixel = 8'hff;
				8'd41:asciipixel = 8'h66;
				8'd42:asciipixel = 8'h65;
				8'd43:asciipixel = 8'hff;
				8'd44:asciipixel = 8'he6;
				8'd45:asciipixel = 8'h25;
				8'd46:asciipixel = 8'h2b;
				8'd47:asciipixel = 8'hea;
				8'd48:asciipixel = 8'h32;
				8'd49:asciipixel = 8'h99;
				8'd50:asciipixel = 8'hff;
				8'd51:asciipixel = 8'h66;
				8'd52:asciipixel = 8'h65;
				8'd53:asciipixel = 8'he9;
				8'd54:asciipixel = 8'h2a;
				8'd55:asciipixel = 8'h26;
				8'd56:asciipixel = 8'he6;
				8'd57:asciipixel = 8'hff;
				8'd58:asciipixel = 8'h32;
				8'd59:asciipixel = 8'h99;
				8'd60:asciipixel = 8'hff;
				8'd61:asciipixel = 8'h74;
				8'd62:asciipixel = 8'h43;
				8'd63:asciipixel = 8'h2e;
				8'd64:asciipixel = 8'h21;
				8'd65:asciipixel = 8'he2;
				8'd66:asciipixel = 8'hff;
				8'd67:asciipixel = 8'hff;
				8'd68:asciipixel = 8'h21;
				8'd69:asciipixel = 8'ha7;
				8'd70:asciipixel = 8'hff;
				8'd71:asciipixel = 8'hb9;
				8'd72:asciipixel = 8'h0;
				8'd73:asciipixel = 8'h10;
				8'd74:asciipixel = 8'hda;
				8'd75:asciipixel = 8'hff;
				8'd76:asciipixel = 8'hf6;
				8'd77:asciipixel = 8'h93;
				8'd78:asciipixel = 8'h6;
				8'd79:asciipixel = 8'he5;
				8'd80:asciipixel = 8'hff;
				8'd81:asciipixel = 8'hfe;
				8'd82:asciipixel = 8'h7a;
				8'd83:asciipixel = 8'h6;
				8'd84:asciipixel = 8'h0;
				8'd85:asciipixel = 8'h0;
				8'd86:asciipixel = 8'h0;
				8'd87:asciipixel = 8'hf;
				8'd88:asciipixel = 8'ha3;
				8'd89:asciipixel = 8'hff;
				8'd90:asciipixel = 8'hff;
				8'd91:asciipixel = 8'hff;
				8'd92:asciipixel = 8'hff;
				8'd93:asciipixel = 8'hf1;
				8'd94:asciipixel = 8'hcf;
				8'd95:asciipixel = 8'hcc;
				8'd96:asciipixel = 8'hd3;
				8'd97:asciipixel = 8'hf8;
				8'd98:asciipixel = 8'hff;
				8'd99:asciipixel = 8'hff;
				default:asciipixel = 0;
			endcase
		end
		else if (num == 'd8) begin // 8
			case(addr)
				8'd00:asciipixel = 8'hff;
				8'd01:asciipixel = 8'hff;
				8'd02:asciipixel = 8'hff;
				8'd03:asciipixel = 8'hff;
				8'd04:asciipixel = 8'hff;
				8'd05:asciipixel = 8'hff;
				8'd06:asciipixel = 8'hff;
				8'd07:asciipixel = 8'hff;
				8'd08:asciipixel = 8'hff;
				8'd09:asciipixel = 8'hff;
				8'd10:asciipixel = 8'hff;
				8'd11:asciipixel = 8'he5;
				8'd12:asciipixel = 8'h32;
				8'd13:asciipixel = 8'h4;
				8'd14:asciipixel = 8'h34;
				8'd15:asciipixel = 8'haf;
				8'd16:asciipixel = 8'h21;
				8'd17:asciipixel = 8'h4;
				8'd18:asciipixel = 8'h4e;
				8'd19:asciipixel = 8'hf9;
				8'd20:asciipixel = 8'hff;
				8'd21:asciipixel = 8'h80;
				8'd22:asciipixel = 8'h2b;
				8'd23:asciipixel = 8'hc2;
				8'd24:asciipixel = 8'h6e;
				8'd25:asciipixel = 8'h8;
				8'd26:asciipixel = 8'h96;
				8'd27:asciipixel = 8'hb7;
				8'd28:asciipixel = 8'he;
				8'd29:asciipixel = 8'hb3;
				8'd30:asciipixel = 8'hff;
				8'd31:asciipixel = 8'h66;
				8'd32:asciipixel = 8'h65;
				8'd33:asciipixel = 8'hff;
				8'd34:asciipixel = 8'hcb;
				8'd35:asciipixel = 8'h0;
				8'd36:asciipixel = 8'hfe;
				8'd37:asciipixel = 8'hff;
				8'd38:asciipixel = 8'h32;
				8'd39:asciipixel = 8'h99;
				8'd40:asciipixel = 8'hff;
				8'd41:asciipixel = 8'h66;
				8'd42:asciipixel = 8'h66;
				8'd43:asciipixel = 8'hff;
				8'd44:asciipixel = 8'hcc;
				8'd45:asciipixel = 8'h0;
				8'd46:asciipixel = 8'hff;
				8'd47:asciipixel = 8'hff;
				8'd48:asciipixel = 8'h33;
				8'd49:asciipixel = 8'h99;
				8'd50:asciipixel = 8'hff;
				8'd51:asciipixel = 8'h66;
				8'd52:asciipixel = 8'h66;
				8'd53:asciipixel = 8'hff;
				8'd54:asciipixel = 8'hcc;
				8'd55:asciipixel = 8'h0;
				8'd56:asciipixel = 8'hff;
				8'd57:asciipixel = 8'hff;
				8'd58:asciipixel = 8'h33;
				8'd59:asciipixel = 8'h99;
				8'd60:asciipixel = 8'hff;
				8'd61:asciipixel = 8'h66;
				8'd62:asciipixel = 8'h66;
				8'd63:asciipixel = 8'hff;
				8'd64:asciipixel = 8'hcb;
				8'd65:asciipixel = 8'h0;
				8'd66:asciipixel = 8'hfe;
				8'd67:asciipixel = 8'hff;
				8'd68:asciipixel = 8'h33;
				8'd69:asciipixel = 8'h99;
				8'd70:asciipixel = 8'hff;
				8'd71:asciipixel = 8'h78;
				8'd72:asciipixel = 8'h3f;
				8'd73:asciipixel = 8'hf5;
				8'd74:asciipixel = 8'h96;
				8'd75:asciipixel = 8'h2;
				8'd76:asciipixel = 8'hc8;
				8'd77:asciipixel = 8'hea;
				8'd78:asciipixel = 8'h18;
				8'd79:asciipixel = 8'ha9;
				8'd80:asciipixel = 8'hff;
				8'd81:asciipixel = 8'hd6;
				8'd82:asciipixel = 8'h13;
				8'd83:asciipixel = 8'h0;
				8'd84:asciipixel = 8'ha;
				8'd85:asciipixel = 8'h80;
				8'd86:asciipixel = 8'h3;
				8'd87:asciipixel = 8'h0;
				8'd88:asciipixel = 8'h22;
				8'd89:asciipixel = 8'hf0;
				8'd90:asciipixel = 8'hff;
				8'd91:asciipixel = 8'hff;
				8'd92:asciipixel = 8'hf4;
				8'd93:asciipixel = 8'hd0;
				8'd94:asciipixel = 8'hee;
				8'd95:asciipixel = 8'hff;
				8'd96:asciipixel = 8'he9;
				8'd97:asciipixel = 8'hd1;
				8'd98:asciipixel = 8'hf8;
				8'd99:asciipixel = 8'hff;
				default:asciipixel = 0;
			endcase
		end
		else if (num == 'd3) begin // 3
			case(addr)
				8'd00:asciipixel = 8'hff;
				8'd01:asciipixel = 8'hef;
				8'd02:asciipixel = 8'hef;
				8'd03:asciipixel = 8'hff;
				8'd04:asciipixel = 8'hff;
				8'd05:asciipixel = 8'hff;
				8'd06:asciipixel = 8'hff;
				8'd07:asciipixel = 8'hff;
				8'd08:asciipixel = 8'hea;
				8'd09:asciipixel = 8'hf4;
				8'd10:asciipixel = 8'hff;
				8'd11:asciipixel = 8'h66;
				8'd12:asciipixel = 8'h66;
				8'd13:asciipixel = 8'hff;
				8'd14:asciipixel = 8'hff;
				8'd15:asciipixel = 8'hff;
				8'd16:asciipixel = 8'hff;
				8'd17:asciipixel = 8'hff;
				8'd18:asciipixel = 8'h33;
				8'd19:asciipixel = 8'h99;
				8'd20:asciipixel = 8'hff;
				8'd21:asciipixel = 8'h66;
				8'd22:asciipixel = 8'h66;
				8'd23:asciipixel = 8'hff;
				8'd24:asciipixel = 8'hcf;
				8'd25:asciipixel = 8'h27;
				8'd26:asciipixel = 8'hff;
				8'd27:asciipixel = 8'hff;
				8'd28:asciipixel = 8'h33;
				8'd29:asciipixel = 8'h99;
				8'd30:asciipixel = 8'hff;
				8'd31:asciipixel = 8'h66;
				8'd32:asciipixel = 8'h66;
				8'd33:asciipixel = 8'hff;
				8'd34:asciipixel = 8'hc6;
				8'd35:asciipixel = 8'h0;
				8'd36:asciipixel = 8'hff;
				8'd37:asciipixel = 8'hff;
				8'd38:asciipixel = 8'h33;
				8'd39:asciipixel = 8'h99;
				8'd40:asciipixel = 8'hff;
				8'd41:asciipixel = 8'h66;
				8'd42:asciipixel = 8'h66;
				8'd43:asciipixel = 8'hff;
				8'd44:asciipixel = 8'hc6;
				8'd45:asciipixel = 8'h0;
				8'd46:asciipixel = 8'hff;
				8'd47:asciipixel = 8'hff;
				8'd48:asciipixel = 8'h33;
				8'd49:asciipixel = 8'h99;
				8'd50:asciipixel = 8'hff;
				8'd51:asciipixel = 8'h66;
				8'd52:asciipixel = 8'h66;
				8'd53:asciipixel = 8'hff;
				8'd54:asciipixel = 8'hc6;
				8'd55:asciipixel = 8'h0;
				8'd56:asciipixel = 8'hff;
				8'd57:asciipixel = 8'hff;
				8'd58:asciipixel = 8'h33;
				8'd59:asciipixel = 8'h99;
				8'd60:asciipixel = 8'hff;
				8'd61:asciipixel = 8'h66;
				8'd62:asciipixel = 8'h65;
				8'd63:asciipixel = 8'hff;
				8'd64:asciipixel = 8'hc5;
				8'd65:asciipixel = 8'h0;
				8'd66:asciipixel = 8'hfe;
				8'd67:asciipixel = 8'hff;
				8'd68:asciipixel = 8'h32;
				8'd69:asciipixel = 8'h99;
				8'd70:asciipixel = 8'hff;
				8'd71:asciipixel = 8'h81;
				8'd72:asciipixel = 8'h2c;
				8'd73:asciipixel = 8'hc3;
				8'd74:asciipixel = 8'h6c;
				8'd75:asciipixel = 8'h8;
				8'd76:asciipixel = 8'h97;
				8'd77:asciipixel = 8'hb8;
				8'd78:asciipixel = 8'hf;
				8'd79:asciipixel = 8'hb2;
				8'd80:asciipixel = 8'hff;
				8'd81:asciipixel = 8'he8;
				8'd82:asciipixel = 8'h3a;
				8'd83:asciipixel = 8'h4;
				8'd84:asciipixel = 8'h2d;
				8'd85:asciipixel = 8'had;
				8'd86:asciipixel = 8'h21;
				8'd87:asciipixel = 8'h5;
				8'd88:asciipixel = 8'h4e;
				8'd89:asciipixel = 8'hf9;
				8'd90:asciipixel = 8'hff;
				8'd91:asciipixel = 8'hff;
				8'd92:asciipixel = 8'hff;
				8'd93:asciipixel = 8'hff;
				8'd94:asciipixel = 8'hff;
				8'd95:asciipixel = 8'hff;
				8'd96:asciipixel = 8'hff;
				8'd97:asciipixel = 8'hff;
				8'd98:asciipixel = 8'hff;
				8'd99:asciipixel = 8'hff;
				default:asciipixel = 0;
			endcase
		end
		else if (num == 'd5) begin // 5
			case(addr)
				8'd00:asciipixel = 8'hff;
				8'd01:asciipixel = 8'hff;
				8'd02:asciipixel = 8'hff;
				8'd03:asciipixel = 8'hff;
				8'd04:asciipixel = 8'hff;
				8'd05:asciipixel = 8'hff;
				8'd06:asciipixel = 8'hff;
				8'd07:asciipixel = 8'hff;
				8'd08:asciipixel = 8'hff;
				8'd09:asciipixel = 8'hff;
				8'd10:asciipixel = 8'hff;
				8'd11:asciipixel = 8'h66;
				8'd12:asciipixel = 8'h0;
				8'd13:asciipixel = 8'h0;
				8'd14:asciipixel = 8'h32;
				8'd15:asciipixel = 8'hff;
				8'd16:asciipixel = 8'hff;
				8'd17:asciipixel = 8'haf;
				8'd18:asciipixel = 8'h70;
				8'd19:asciipixel = 8'hff;
				8'd20:asciipixel = 8'hff;
				8'd21:asciipixel = 8'h66;
				8'd22:asciipixel = 8'h51;
				8'd23:asciipixel = 8'had;
				8'd24:asciipixel = 8'h22;
				8'd25:asciipixel = 8'hff;
				8'd26:asciipixel = 8'hff;
				8'd27:asciipixel = 8'hbb;
				8'd28:asciipixel = 8'h4;
				8'd29:asciipixel = 8'hec;
				8'd30:asciipixel = 8'hff;
				8'd31:asciipixel = 8'h66;
				8'd32:asciipixel = 8'h66;
				8'd33:asciipixel = 8'hdf;
				8'd34:asciipixel = 8'hd;
				8'd35:asciipixel = 8'hff;
				8'd36:asciipixel = 8'hff;
				8'd37:asciipixel = 8'hfe;
				8'd38:asciipixel = 8'h13;
				8'd39:asciipixel = 8'hb5;
				8'd40:asciipixel = 8'hff;
				8'd41:asciipixel = 8'h66;
				8'd42:asciipixel = 8'h66;
				8'd43:asciipixel = 8'hf0;
				8'd44:asciipixel = 8'h0;
				8'd45:asciipixel = 8'hef;
				8'd46:asciipixel = 8'hff;
				8'd47:asciipixel = 8'hff;
				8'd48:asciipixel = 8'h2e;
				8'd49:asciipixel = 8'h9d;
				8'd50:asciipixel = 8'hff;
				8'd51:asciipixel = 8'h66;
				8'd52:asciipixel = 8'h66;
				8'd53:asciipixel = 8'hfe;
				8'd54:asciipixel = 8'h10;
				8'd55:asciipixel = 8'hc6;
				8'd56:asciipixel = 8'hff;
				8'd57:asciipixel = 8'hff;
				8'd58:asciipixel = 8'h2d;
				8'd59:asciipixel = 8'h9c;
				8'd60:asciipixel = 8'hff;
				8'd61:asciipixel = 8'h66;
				8'd62:asciipixel = 8'h66;
				8'd63:asciipixel = 8'hff;
				8'd64:asciipixel = 8'h44;
				8'd65:asciipixel = 8'h89;
				8'd66:asciipixel = 8'hff;
				8'd67:asciipixel = 8'hf5;
				8'd68:asciipixel = 8'ha;
				8'd69:asciipixel = 8'hb7;
				8'd70:asciipixel = 8'hff;
				8'd71:asciipixel = 8'h66;
				8'd72:asciipixel = 8'h66;
				8'd73:asciipixel = 8'hff;
				8'd74:asciipixel = 8'h9a;
				8'd75:asciipixel = 8'h20;
				8'd76:asciipixel = 8'hd0;
				8'd77:asciipixel = 8'h60;
				8'd78:asciipixel = 8'hd;
				8'd79:asciipixel = 8'hf1;
				8'd80:asciipixel = 8'hff;
				8'd81:asciipixel = 8'h66;
				8'd82:asciipixel = 8'h66;
				8'd83:asciipixel = 8'hff;
				8'd84:asciipixel = 8'hfa;
				8'd85:asciipixel = 8'h4e;
				8'd86:asciipixel = 8'h0;
				8'd87:asciipixel = 8'hf;
				8'd88:asciipixel = 8'haa;
				8'd89:asciipixel = 8'hff;
				8'd90:asciipixel = 8'hff;
				8'd91:asciipixel = 8'hef;
				8'd92:asciipixel = 8'hef;
				8'd93:asciipixel = 8'hff;
				8'd94:asciipixel = 8'hff;
				8'd95:asciipixel = 8'hff;
				8'd96:asciipixel = 8'hec;
				8'd97:asciipixel = 8'hfa;
				8'd98:asciipixel = 8'hff;
				8'd99:asciipixel = 8'hff;
				default:asciipixel = 0;
			endcase
		end
		else if (num == 'd6) begin // 6
			case(addr)
				8'd00:asciipixel = 8'hff;
				8'd01:asciipixel = 8'hff;
				8'd02:asciipixel = 8'hff;
				8'd03:asciipixel = 8'hff;
				8'd04:asciipixel = 8'hff;
				8'd05:asciipixel = 8'hff;
				8'd06:asciipixel = 8'hff;
				8'd07:asciipixel = 8'hff;
				8'd08:asciipixel = 8'hff;
				8'd09:asciipixel = 8'hff;
				8'd10:asciipixel = 8'hff;
				8'd11:asciipixel = 8'hff;
				8'd12:asciipixel = 8'hf6;
				8'd13:asciipixel = 8'h72;
				8'd14:asciipixel = 8'h18;
				8'd15:asciipixel = 8'h1;
				8'd16:asciipixel = 8'hd;
				8'd17:asciipixel = 8'h39;
				8'd18:asciipixel = 8'ha3;
				8'd19:asciipixel = 8'hff;
				8'd20:asciipixel = 8'hff;
				8'd21:asciipixel = 8'hff;
				8'd22:asciipixel = 8'h5a;
				8'd23:asciipixel = 8'h24;
				8'd24:asciipixel = 8'h73;
				8'd25:asciipixel = 8'h0;
				8'd26:asciipixel = 8'h6f;
				8'd27:asciipixel = 8'h50;
				8'd28:asciipixel = 8'h0;
				8'd29:asciipixel = 8'hc0;
				8'd30:asciipixel = 8'hff;
				8'd31:asciipixel = 8'hd9;
				8'd32:asciipixel = 8'h1;
				8'd33:asciipixel = 8'hce;
				8'd34:asciipixel = 8'hcb;
				8'd35:asciipixel = 8'h0;
				8'd36:asciipixel = 8'hfe;
				8'd37:asciipixel = 8'hff;
				8'd38:asciipixel = 8'h2f;
				8'd39:asciipixel = 8'h99;
				8'd40:asciipixel = 8'hff;
				8'd41:asciipixel = 8'h94;
				8'd42:asciipixel = 8'h2d;
				8'd43:asciipixel = 8'hff;
				8'd44:asciipixel = 8'hcc;
				8'd45:asciipixel = 8'h0;
				8'd46:asciipixel = 8'hff;
				8'd47:asciipixel = 8'hff;
				8'd48:asciipixel = 8'h33;
				8'd49:asciipixel = 8'h99;
				8'd50:asciipixel = 8'hff;
				8'd51:asciipixel = 8'h72;
				8'd52:asciipixel = 8'h57;
				8'd53:asciipixel = 8'hff;
				8'd54:asciipixel = 8'hcc;
				8'd55:asciipixel = 8'h0;
				8'd56:asciipixel = 8'hff;
				8'd57:asciipixel = 8'hff;
				8'd58:asciipixel = 8'h33;
				8'd59:asciipixel = 8'h99;
				8'd60:asciipixel = 8'hff;
				8'd61:asciipixel = 8'ha4;
				8'd62:asciipixel = 8'ha1;
				8'd63:asciipixel = 8'hff;
				8'd64:asciipixel = 8'hcc;
				8'd65:asciipixel = 8'h0;
				8'd66:asciipixel = 8'hff;
				8'd67:asciipixel = 8'hff;
				8'd68:asciipixel = 8'h33;
				8'd69:asciipixel = 8'h99;
				8'd70:asciipixel = 8'hff;
				8'd71:asciipixel = 8'hff;
				8'd72:asciipixel = 8'hff;
				8'd73:asciipixel = 8'hff;
				8'd74:asciipixel = 8'hdc;
				8'd75:asciipixel = 8'h0;
				8'd76:asciipixel = 8'hd1;
				8'd77:asciipixel = 8'heb;
				8'd78:asciipixel = 8'h19;
				8'd79:asciipixel = 8'ha7;
				8'd80:asciipixel = 8'hff;
				8'd81:asciipixel = 8'hff;
				8'd82:asciipixel = 8'hff;
				8'd83:asciipixel = 8'hff;
				8'd84:asciipixel = 8'hfe;
				8'd85:asciipixel = 8'h54;
				8'd86:asciipixel = 8'h0;
				8'd87:asciipixel = 8'h0;
				8'd88:asciipixel = 8'h2b;
				8'd89:asciipixel = 8'hf0;
				8'd90:asciipixel = 8'hff;
				8'd91:asciipixel = 8'hff;
				8'd92:asciipixel = 8'hff;
				8'd93:asciipixel = 8'hff;
				8'd94:asciipixel = 8'hff;
				8'd95:asciipixel = 8'hfe;
				8'd96:asciipixel = 8'hdc;
				8'd97:asciipixel = 8'hd5;
				8'd98:asciipixel = 8'hfb;
				8'd99:asciipixel = 8'hff;
				default:asciipixel = 0;
			endcase
		end
		else if (num == 'd9) begin // 9
			case(addr)
				8'd00:asciipixel = 8'hff;
				8'd01:asciipixel = 8'hff;
				8'd02:asciipixel = 8'hff;
				8'd03:asciipixel = 8'hff;
				8'd04:asciipixel = 8'hff;
				8'd05:asciipixel = 8'hff;
				8'd06:asciipixel = 8'hff;
				8'd07:asciipixel = 8'hff;
				8'd08:asciipixel = 8'hff;
				8'd09:asciipixel = 8'hff;
				8'd10:asciipixel = 8'hff;
				8'd11:asciipixel = 8'he8;
				8'd12:asciipixel = 8'h3e;
				8'd13:asciipixel = 8'h5;
				8'd14:asciipixel = 8'h1b;
				8'd15:asciipixel = 8'hac;
				8'd16:asciipixel = 8'hff;
				8'd17:asciipixel = 8'hff;
				8'd18:asciipixel = 8'hff;
				8'd19:asciipixel = 8'hff;
				8'd20:asciipixel = 8'hff;
				8'd21:asciipixel = 8'h7e;
				8'd22:asciipixel = 8'h2c;
				8'd23:asciipixel = 8'hc3;
				8'd24:asciipixel = 8'h77;
				8'd25:asciipixel = 8'h1b;
				8'd26:asciipixel = 8'hff;
				8'd27:asciipixel = 8'hff;
				8'd28:asciipixel = 8'hff;
				8'd29:asciipixel = 8'hff;
				8'd30:asciipixel = 8'hff;
				8'd31:asciipixel = 8'h66;
				8'd32:asciipixel = 8'h65;
				8'd33:asciipixel = 8'hff;
				8'd34:asciipixel = 8'hcb;
				8'd35:asciipixel = 8'h0;
				8'd36:asciipixel = 8'hff;
				8'd37:asciipixel = 8'hff;
				8'd38:asciipixel = 8'hac;
				8'd39:asciipixel = 8'hd6;
				8'd40:asciipixel = 8'hff;
				8'd41:asciipixel = 8'h66;
				8'd42:asciipixel = 8'h66;
				8'd43:asciipixel = 8'hff;
				8'd44:asciipixel = 8'hcc;
				8'd45:asciipixel = 8'h0;
				8'd46:asciipixel = 8'hff;
				8'd47:asciipixel = 8'hff;
				8'd48:asciipixel = 8'h29;
				8'd49:asciipixel = 8'ha1;
				8'd50:asciipixel = 8'hff;
				8'd51:asciipixel = 8'h66;
				8'd52:asciipixel = 8'h66;
				8'd53:asciipixel = 8'hff;
				8'd54:asciipixel = 8'hcc;
				8'd55:asciipixel = 8'h0;
				8'd56:asciipixel = 8'hff;
				8'd57:asciipixel = 8'hfb;
				8'd58:asciipixel = 8'ha;
				8'd59:asciipixel = 8'hbe;
				8'd60:asciipixel = 8'hff;
				8'd61:asciipixel = 8'h66;
				8'd62:asciipixel = 8'h65;
				8'd63:asciipixel = 8'hff;
				8'd64:asciipixel = 8'hcb;
				8'd65:asciipixel = 8'h0;
				8'd66:asciipixel = 8'hff;
				8'd67:asciipixel = 8'hb5;
				8'd68:asciipixel = 8'h8;
				8'd69:asciipixel = 8'hf2;
				8'd70:asciipixel = 8'hff;
				8'd71:asciipixel = 8'h7c;
				8'd72:asciipixel = 8'h17;
				8'd73:asciipixel = 8'h96;
				8'd74:asciipixel = 8'h7d;
				8'd75:asciipixel = 8'h0;
				8'd76:asciipixel = 8'hba;
				8'd77:asciipixel = 8'h22;
				8'd78:asciipixel = 8'h6c;
				8'd79:asciipixel = 8'hff;
				8'd80:asciipixel = 8'hff;
				8'd81:asciipixel = 8'hee;
				8'd82:asciipixel = 8'h52;
				8'd83:asciipixel = 8'h4;
				8'd84:asciipixel = 8'h0;
				8'd85:asciipixel = 8'h0;
				8'd86:asciipixel = 8'h2;
				8'd87:asciipixel = 8'h5e;
				8'd88:asciipixel = 8'hf6;
				8'd89:asciipixel = 8'hff;
				8'd90:asciipixel = 8'hff;
				8'd91:asciipixel = 8'hff;
				8'd92:asciipixel = 8'hff;
				8'd93:asciipixel = 8'hf4;
				8'd94:asciipixel = 8'hd5;
				8'd95:asciipixel = 8'hce;
				8'd96:asciipixel = 8'hed;
				8'd97:asciipixel = 8'hff;
				8'd98:asciipixel = 8'hff;
				8'd99:asciipixel = 8'hff;
				default:asciipixel = 0;
			endcase
		end
		else if (num == 'd2) begin // 2
			case(addr)
				8'd00:asciipixel = 8'hff;
				8'd01:asciipixel = 8'hff;
				8'd02:asciipixel = 8'hff;
				8'd03:asciipixel = 8'hff;
				8'd04:asciipixel = 8'hff;
				8'd05:asciipixel = 8'hff;
				8'd06:asciipixel = 8'hff;
				8'd07:asciipixel = 8'hff;
				8'd08:asciipixel = 8'hff;
				8'd09:asciipixel = 8'hff;
				8'd10:asciipixel = 8'hff;
				8'd11:asciipixel = 8'hfd;
				8'd12:asciipixel = 8'h4e;
				8'd13:asciipixel = 8'hd2;
				8'd14:asciipixel = 8'hff;
				8'd15:asciipixel = 8'hff;
				8'd16:asciipixel = 8'hff;
				8'd17:asciipixel = 8'h88;
				8'd18:asciipixel = 8'h0;
				8'd19:asciipixel = 8'h99;
				8'd20:asciipixel = 8'hff;
				8'd21:asciipixel = 8'hbf;
				8'd22:asciipixel = 8'h9;
				8'd23:asciipixel = 8'he4;
				8'd24:asciipixel = 8'hff;
				8'd25:asciipixel = 8'hff;
				8'd26:asciipixel = 8'hfd;
				8'd27:asciipixel = 8'h23;
				8'd28:asciipixel = 8'h0;
				8'd29:asciipixel = 8'h99;
				8'd30:asciipixel = 8'hff;
				8'd31:asciipixel = 8'h84;
				8'd32:asciipixel = 8'h45;
				8'd33:asciipixel = 8'hff;
				8'd34:asciipixel = 8'hff;
				8'd35:asciipixel = 8'hff;
				8'd36:asciipixel = 8'hb5;
				8'd37:asciipixel = 8'h10;
				8'd38:asciipixel = 8'h2a;
				8'd39:asciipixel = 8'h99;
				8'd40:asciipixel = 8'hff;
				8'd41:asciipixel = 8'h6b;
				8'd42:asciipixel = 8'h61;
				8'd43:asciipixel = 8'hff;
				8'd44:asciipixel = 8'hff;
				8'd45:asciipixel = 8'hff;
				8'd46:asciipixel = 8'h43;
				8'd47:asciipixel = 8'h6c;
				8'd48:asciipixel = 8'h33;
				8'd49:asciipixel = 8'h99;
				8'd50:asciipixel = 8'hff;
				8'd51:asciipixel = 8'h69;
				8'd52:asciipixel = 8'h61;
				8'd53:asciipixel = 8'hff;
				8'd54:asciipixel = 8'hff;
				8'd55:asciipixel = 8'hc6;
				8'd56:asciipixel = 8'h2;
				8'd57:asciipixel = 8'hd7;
				8'd58:asciipixel = 8'h33;
				8'd59:asciipixel = 8'h99;
				8'd60:asciipixel = 8'hff;
				8'd61:asciipixel = 8'h81;
				8'd62:asciipixel = 8'h3f;
				8'd63:asciipixel = 8'hff;
				8'd64:asciipixel = 8'hfd;
				8'd65:asciipixel = 8'h3a;
				8'd66:asciipixel = 8'h55;
				8'd67:asciipixel = 8'hff;
				8'd68:asciipixel = 8'h33;
				8'd69:asciipixel = 8'h99;
				8'd70:asciipixel = 8'hff;
				8'd71:asciipixel = 8'hc4;
				8'd72:asciipixel = 8'h3;
				8'd73:asciipixel = 8'hb0;
				8'd74:asciipixel = 8'h77;
				8'd75:asciipixel = 8'h8;
				8'd76:asciipixel = 8'hdb;
				8'd77:asciipixel = 8'hff;
				8'd78:asciipixel = 8'h33;
				8'd79:asciipixel = 8'h99;
				8'd80:asciipixel = 8'hff;
				8'd81:asciipixel = 8'hff;
				8'd82:asciipixel = 8'h6a;
				8'd83:asciipixel = 8'h0;
				8'd84:asciipixel = 8'h3;
				8'd85:asciipixel = 8'ha1;
				8'd86:asciipixel = 8'hff;
				8'd87:asciipixel = 8'hff;
				8'd88:asciipixel = 8'h33;
				8'd89:asciipixel = 8'h99;
				8'd90:asciipixel = 8'hff;
				8'd91:asciipixel = 8'hff;
				8'd92:asciipixel = 8'hff;
				8'd93:asciipixel = 8'he2;
				8'd94:asciipixel = 8'he1;
				8'd95:asciipixel = 8'hff;
				8'd96:asciipixel = 8'hff;
				8'd97:asciipixel = 8'hff;
				8'd98:asciipixel = 8'hd6;
				8'd99:asciipixel = 8'hea;
				default:asciipixel = 0;
			endcase
		end
		else if (num == 'd4) begin // 4
			case(addr)
				8'd00:asciipixel = 8'hff;
				8'd01:asciipixel = 8'hff;
				8'd02:asciipixel = 8'hff;
				8'd03:asciipixel = 8'hff;
				8'd04:asciipixel = 8'hff;
				8'd05:asciipixel = 8'hff;
				8'd06:asciipixel = 8'hff;
				8'd07:asciipixel = 8'hff;
				8'd08:asciipixel = 8'hff;
				8'd09:asciipixel = 8'hff;
				8'd10:asciipixel = 8'hff;
				8'd11:asciipixel = 8'hff;
				8'd12:asciipixel = 8'hff;
				8'd13:asciipixel = 8'hff;
				8'd14:asciipixel = 8'hdd;
				8'd15:asciipixel = 8'hf;
				8'd16:asciipixel = 8'h33;
				8'd17:asciipixel = 8'hff;
				8'd18:asciipixel = 8'hff;
				8'd19:asciipixel = 8'hff;
				8'd20:asciipixel = 8'hff;
				8'd21:asciipixel = 8'hff;
				8'd22:asciipixel = 8'hff;
				8'd23:asciipixel = 8'hf9;
				8'd24:asciipixel = 8'h36;
				8'd25:asciipixel = 8'h10;
				8'd26:asciipixel = 8'h33;
				8'd27:asciipixel = 8'hff;
				8'd28:asciipixel = 8'hff;
				8'd29:asciipixel = 8'hff;
				8'd30:asciipixel = 8'hff;
				8'd31:asciipixel = 8'hff;
				8'd32:asciipixel = 8'hff;
				8'd33:asciipixel = 8'h74;
				8'd34:asciipixel = 8'h19;
				8'd35:asciipixel = 8'h87;
				8'd36:asciipixel = 8'h33;
				8'd37:asciipixel = 8'hff;
				8'd38:asciipixel = 8'hff;
				8'd39:asciipixel = 8'hff;
				8'd40:asciipixel = 8'hff;
				8'd41:asciipixel = 8'hff;
				8'd42:asciipixel = 8'hb6;
				8'd43:asciipixel = 8'h1;
				8'd44:asciipixel = 8'hb1;
				8'd45:asciipixel = 8'h99;
				8'd46:asciipixel = 8'h33;
				8'd47:asciipixel = 8'hff;
				8'd48:asciipixel = 8'hff;
				8'd49:asciipixel = 8'hff;
				8'd50:asciipixel = 8'hff;
				8'd51:asciipixel = 8'he5;
				8'd52:asciipixel = 8'h15;
				8'd53:asciipixel = 8'h5d;
				8'd54:asciipixel = 8'hff;
				8'd55:asciipixel = 8'h99;
				8'd56:asciipixel = 8'h33;
				8'd57:asciipixel = 8'hff;
				8'd58:asciipixel = 8'hff;
				8'd59:asciipixel = 8'hff;
				8'd60:asciipixel = 8'hff;
				8'd61:asciipixel = 8'h6d;
				8'd62:asciipixel = 8'h1;
				8'd63:asciipixel = 8'h87;
				8'd64:asciipixel = 8'h99;
				8'd65:asciipixel = 8'h5b;
				8'd66:asciipixel = 8'h1e;
				8'd67:asciipixel = 8'h99;
				8'd68:asciipixel = 8'h99;
				8'd69:asciipixel = 8'hd6;
				8'd70:asciipixel = 8'hff;
				8'd71:asciipixel = 8'h84;
				8'd72:asciipixel = 8'h33;
				8'd73:asciipixel = 8'h33;
				8'd74:asciipixel = 8'h33;
				8'd75:asciipixel = 8'h1e;
				8'd76:asciipixel = 8'ha;
				8'd77:asciipixel = 8'h33;
				8'd78:asciipixel = 8'h33;
				8'd79:asciipixel = 8'had;
				8'd80:asciipixel = 8'hff;
				8'd81:asciipixel = 8'hff;
				8'd82:asciipixel = 8'hff;
				8'd83:asciipixel = 8'hff;
				8'd84:asciipixel = 8'hff;
				8'd85:asciipixel = 8'h99;
				8'd86:asciipixel = 8'h33;
				8'd87:asciipixel = 8'hff;
				8'd88:asciipixel = 8'hff;
				8'd89:asciipixel = 8'hff;
				8'd90:asciipixel = 8'hff;
				8'd91:asciipixel = 8'hff;
				8'd92:asciipixel = 8'hff;
				8'd93:asciipixel = 8'hff;
				8'd94:asciipixel = 8'hff;
				8'd95:asciipixel = 8'hf4;
				8'd96:asciipixel = 8'hea;
				8'd97:asciipixel = 8'hff;
				8'd98:asciipixel = 8'hff;
				8'd99:asciipixel = 8'hff;
				default:asciipixel = 0;
			endcase
		end
		else if (num == 'd13) begin // *
			case(addr)
				8'd00:asciipixel = 8'hff;
				8'd01:asciipixel = 8'hff;
				8'd02:asciipixel = 8'hff;
				8'd03:asciipixel = 8'hff;
				8'd04:asciipixel = 8'hff;
				8'd05:asciipixel = 8'hff;
				8'd06:asciipixel = 8'hff;
				8'd07:asciipixel = 8'hff;
				8'd08:asciipixel = 8'hff;
				8'd09:asciipixel = 8'hff;
				8'd10:asciipixel = 8'hff;
				8'd11:asciipixel = 8'hff;
				8'd12:asciipixel = 8'hfe;
				8'd13:asciipixel = 8'hff;
				8'd14:asciipixel = 8'hcc;
				8'd15:asciipixel = 8'h0;
				8'd16:asciipixel = 8'hff;
				8'd17:asciipixel = 8'hfe;
				8'd18:asciipixel = 8'hff;
				8'd19:asciipixel = 8'hff;
				8'd20:asciipixel = 8'hff;
				8'd21:asciipixel = 8'hff;
				8'd22:asciipixel = 8'h68;
				8'd23:asciipixel = 8'h6b;
				8'd24:asciipixel = 8'hc8;
				8'd25:asciipixel = 8'h0;
				8'd26:asciipixel = 8'hee;
				8'd27:asciipixel = 8'h45;
				8'd28:asciipixel = 8'h99;
				8'd29:asciipixel = 8'hff;
				8'd30:asciipixel = 8'hff;
				8'd31:asciipixel = 8'hff;
				8'd32:asciipixel = 8'hb5;
				8'd33:asciipixel = 8'h10;
				8'd34:asciipixel = 8'h29;
				8'd35:asciipixel = 8'h0;
				8'd36:asciipixel = 8'h27;
				8'd37:asciipixel = 8'h25;
				8'd38:asciipixel = 8'hd3;
				8'd39:asciipixel = 8'hff;
				8'd40:asciipixel = 8'hff;
				8'd41:asciipixel = 8'hff;
				8'd42:asciipixel = 8'hff;
				8'd43:asciipixel = 8'hdb;
				8'd44:asciipixel = 8'h2d;
				8'd45:asciipixel = 8'h0;
				8'd46:asciipixel = 8'h4c;
				8'd47:asciipixel = 8'hef;
				8'd48:asciipixel = 8'hff;
				8'd49:asciipixel = 8'hff;
				8'd50:asciipixel = 8'hff;
				8'd51:asciipixel = 8'hff;
				8'd52:asciipixel = 8'hff;
				8'd53:asciipixel = 8'hf3;
				8'd54:asciipixel = 8'h53;
				8'd55:asciipixel = 8'h0;
				8'd56:asciipixel = 8'h7c;
				8'd57:asciipixel = 8'hfd;
				8'd58:asciipixel = 8'hff;
				8'd59:asciipixel = 8'hff;
				8'd60:asciipixel = 8'hff;
				8'd61:asciipixel = 8'hff;
				8'd62:asciipixel = 8'hda;
				8'd63:asciipixel = 8'h2c;
				8'd64:asciipixel = 8'hf;
				8'd65:asciipixel = 8'h0;
				8'd66:asciipixel = 8'hf;
				8'd67:asciipixel = 8'h4a;
				8'd68:asciipixel = 8'hee;
				8'd69:asciipixel = 8'hff;
				8'd70:asciipixel = 8'hff;
				8'd71:asciipixel = 8'hff;
				8'd72:asciipixel = 8'h4d;
				8'd73:asciipixel = 8'h3e;
				8'd74:asciipixel = 8'hb9;
				8'd75:asciipixel = 8'h0;
				8'd76:asciipixel = 8'hd5;
				8'd77:asciipixel = 8'h22;
				8'd78:asciipixel = 8'h80;
				8'd79:asciipixel = 8'hff;
				8'd80:asciipixel = 8'hff;
				8'd81:asciipixel = 8'hff;
				8'd82:asciipixel = 8'hf3;
				8'd83:asciipixel = 8'hf9;
				8'd84:asciipixel = 8'hcc;
				8'd85:asciipixel = 8'h0;
				8'd86:asciipixel = 8'hff;
				8'd87:asciipixel = 8'hee;
				8'd88:asciipixel = 8'hfd;
				8'd89:asciipixel = 8'hff;
				8'd90:asciipixel = 8'hff;
				8'd91:asciipixel = 8'hff;
				8'd92:asciipixel = 8'hff;
				8'd93:asciipixel = 8'hff;
				8'd94:asciipixel = 8'hf4;
				8'd95:asciipixel = 8'hcc;
				8'd96:asciipixel = 8'hff;
				8'd97:asciipixel = 8'hff;
				8'd98:asciipixel = 8'hff;
				8'd99:asciipixel = 8'hff;
				default:asciipixel = 0;
			endcase
		end
		else if (num == 'd1) begin // 1
			case(addr)
				8'd00:asciipixel = 8'hff;
				8'd01:asciipixel = 8'hff;
				8'd02:asciipixel = 8'hff;
				8'd03:asciipixel = 8'hff;
				8'd04:asciipixel = 8'hff;
				8'd05:asciipixel = 8'hff;
				8'd06:asciipixel = 8'hff;
				8'd07:asciipixel = 8'hff;
				8'd08:asciipixel = 8'hff;
				8'd09:asciipixel = 8'hff;
				8'd10:asciipixel = 8'hff;
				8'd11:asciipixel = 8'hff;
				8'd12:asciipixel = 8'hff;
				8'd13:asciipixel = 8'hff;
				8'd14:asciipixel = 8'hff;
				8'd15:asciipixel = 8'hff;
				8'd16:asciipixel = 8'hff;
				8'd17:asciipixel = 8'hff;
				8'd18:asciipixel = 8'h33;
				8'd19:asciipixel = 8'h99;
				8'd20:asciipixel = 8'hff;
				8'd21:asciipixel = 8'hff;
				8'd22:asciipixel = 8'hef;
				8'd23:asciipixel = 8'hd9;
				8'd24:asciipixel = 8'hfa;
				8'd25:asciipixel = 8'hff;
				8'd26:asciipixel = 8'hff;
				8'd27:asciipixel = 8'hff;
				8'd28:asciipixel = 8'h33;
				8'd29:asciipixel = 8'h99;
				8'd30:asciipixel = 8'hff;
				8'd31:asciipixel = 8'hf2;
				8'd32:asciipixel = 8'h2b;
				8'd33:asciipixel = 8'h56;
				8'd34:asciipixel = 8'hfe;
				8'd35:asciipixel = 8'hff;
				8'd36:asciipixel = 8'hff;
				8'd37:asciipixel = 8'hff;
				8'd38:asciipixel = 8'h33;
				8'd39:asciipixel = 8'h99;
				8'd40:asciipixel = 8'hff;
				8'd41:asciipixel = 8'h76;
				8'd42:asciipixel = 8'h0;
				8'd43:asciipixel = 8'h5a;
				8'd44:asciipixel = 8'h66;
				8'd45:asciipixel = 8'h66;
				8'd46:asciipixel = 8'h66;
				8'd47:asciipixel = 8'h66;
				8'd48:asciipixel = 8'h14;
				8'd49:asciipixel = 8'h99;
				8'd50:asciipixel = 8'hff;
				8'd51:asciipixel = 8'ha3;
				8'd52:asciipixel = 8'h66;
				8'd53:asciipixel = 8'h66;
				8'd54:asciipixel = 8'h66;
				8'd55:asciipixel = 8'h66;
				8'd56:asciipixel = 8'h66;
				8'd57:asciipixel = 8'h66;
				8'd58:asciipixel = 8'h14;
				8'd59:asciipixel = 8'h99;
				8'd60:asciipixel = 8'hff;
				8'd61:asciipixel = 8'hff;
				8'd62:asciipixel = 8'hff;
				8'd63:asciipixel = 8'hff;
				8'd64:asciipixel = 8'hff;
				8'd65:asciipixel = 8'hff;
				8'd66:asciipixel = 8'hff;
				8'd67:asciipixel = 8'hff;
				8'd68:asciipixel = 8'h33;
				8'd69:asciipixel = 8'h99;
				8'd70:asciipixel = 8'hff;
				8'd71:asciipixel = 8'hff;
				8'd72:asciipixel = 8'hff;
				8'd73:asciipixel = 8'hff;
				8'd74:asciipixel = 8'hff;
				8'd75:asciipixel = 8'hff;
				8'd76:asciipixel = 8'hff;
				8'd77:asciipixel = 8'hff;
				8'd78:asciipixel = 8'h33;
				8'd79:asciipixel = 8'h99;
				8'd80:asciipixel = 8'hff;
				8'd81:asciipixel = 8'hff;
				8'd82:asciipixel = 8'hff;
				8'd83:asciipixel = 8'hff;
				8'd84:asciipixel = 8'hff;
				8'd85:asciipixel = 8'hff;
				8'd86:asciipixel = 8'hff;
				8'd87:asciipixel = 8'hff;
				8'd88:asciipixel = 8'h33;
				8'd89:asciipixel = 8'h99;
				8'd90:asciipixel = 8'hff;
				8'd91:asciipixel = 8'hff;
				8'd92:asciipixel = 8'hff;
				8'd93:asciipixel = 8'hff;
				8'd94:asciipixel = 8'hff;
				8'd95:asciipixel = 8'hff;
				8'd96:asciipixel = 8'hff;
				8'd97:asciipixel = 8'hff;
				8'd98:asciipixel = 8'hd6;
				8'd99:asciipixel = 8'hea;
				default:asciipixel = 0;
			endcase
		end
		else if (num == 'd10) begin // =
			case(addr)
				8'd00:asciipixel = 8'hff;
				8'd01:asciipixel = 8'hff;
				8'd02:asciipixel = 8'hff;
				8'd03:asciipixel = 8'hff;
				8'd04:asciipixel = 8'hff;
				8'd05:asciipixel = 8'hff;
				8'd06:asciipixel = 8'hff;
				8'd07:asciipixel = 8'hff;
				8'd08:asciipixel = 8'hff;
				8'd09:asciipixel = 8'hff;
				8'd10:asciipixel = 8'hff;
				8'd11:asciipixel = 8'hff;
				8'd12:asciipixel = 8'hcc;
				8'd13:asciipixel = 8'h0;
				8'd14:asciipixel = 8'hff;
				8'd15:asciipixel = 8'hff;
				8'd16:asciipixel = 8'h99;
				8'd17:asciipixel = 8'h33;
				8'd18:asciipixel = 8'hff;
				8'd19:asciipixel = 8'hff;
				8'd20:asciipixel = 8'hff;
				8'd21:asciipixel = 8'hff;
				8'd22:asciipixel = 8'hcc;
				8'd23:asciipixel = 8'h0;
				8'd24:asciipixel = 8'hff;
				8'd25:asciipixel = 8'hff;
				8'd26:asciipixel = 8'h99;
				8'd27:asciipixel = 8'h33;
				8'd28:asciipixel = 8'hff;
				8'd29:asciipixel = 8'hff;
				8'd30:asciipixel = 8'hff;
				8'd31:asciipixel = 8'hff;
				8'd32:asciipixel = 8'hcc;
				8'd33:asciipixel = 8'h0;
				8'd34:asciipixel = 8'hff;
				8'd35:asciipixel = 8'hff;
				8'd36:asciipixel = 8'h99;
				8'd37:asciipixel = 8'h33;
				8'd38:asciipixel = 8'hff;
				8'd39:asciipixel = 8'hff;
				8'd40:asciipixel = 8'hff;
				8'd41:asciipixel = 8'hff;
				8'd42:asciipixel = 8'hcc;
				8'd43:asciipixel = 8'h0;
				8'd44:asciipixel = 8'hff;
				8'd45:asciipixel = 8'hff;
				8'd46:asciipixel = 8'h99;
				8'd47:asciipixel = 8'h33;
				8'd48:asciipixel = 8'hff;
				8'd49:asciipixel = 8'hff;
				8'd50:asciipixel = 8'hff;
				8'd51:asciipixel = 8'hff;
				8'd52:asciipixel = 8'hcc;
				8'd53:asciipixel = 8'h0;
				8'd54:asciipixel = 8'hff;
				8'd55:asciipixel = 8'hff;
				8'd56:asciipixel = 8'h99;
				8'd57:asciipixel = 8'h33;
				8'd58:asciipixel = 8'hff;
				8'd59:asciipixel = 8'hff;
				8'd60:asciipixel = 8'hff;
				8'd61:asciipixel = 8'hff;
				8'd62:asciipixel = 8'hcc;
				8'd63:asciipixel = 8'h0;
				8'd64:asciipixel = 8'hff;
				8'd65:asciipixel = 8'hff;
				8'd66:asciipixel = 8'h99;
				8'd67:asciipixel = 8'h33;
				8'd68:asciipixel = 8'hff;
				8'd69:asciipixel = 8'hff;
				8'd70:asciipixel = 8'hff;
				8'd71:asciipixel = 8'hff;
				8'd72:asciipixel = 8'hcc;
				8'd73:asciipixel = 8'h0;
				8'd74:asciipixel = 8'hff;
				8'd75:asciipixel = 8'hff;
				8'd76:asciipixel = 8'h99;
				8'd77:asciipixel = 8'h33;
				8'd78:asciipixel = 8'hff;
				8'd79:asciipixel = 8'hff;
				8'd80:asciipixel = 8'hff;
				8'd81:asciipixel = 8'hff;
				8'd82:asciipixel = 8'hcc;
				8'd83:asciipixel = 8'h0;
				8'd84:asciipixel = 8'hff;
				8'd85:asciipixel = 8'hff;
				8'd86:asciipixel = 8'h99;
				8'd87:asciipixel = 8'h33;
				8'd88:asciipixel = 8'hff;
				8'd89:asciipixel = 8'hff;
				8'd90:asciipixel = 8'hff;
				8'd91:asciipixel = 8'hff;
				8'd92:asciipixel = 8'hf4;
				8'd93:asciipixel = 8'hcc;
				8'd94:asciipixel = 8'hff;
				8'd95:asciipixel = 8'hff;
				8'd96:asciipixel = 8'hea;
				8'd97:asciipixel = 8'hd6;
				8'd98:asciipixel = 8'hff;
				8'd99:asciipixel = 8'hff;
				default:asciipixel = 0;
			endcase
		end
		else if (num == 'd7) begin // 7
			case(addr)
				8'd00:asciipixel = 8'hff;
				8'd01:asciipixel = 8'hff;
				8'd02:asciipixel = 8'hff;
				8'd03:asciipixel = 8'hff;
				8'd04:asciipixel = 8'hff;
				8'd05:asciipixel = 8'hff;
				8'd06:asciipixel = 8'hff;
				8'd07:asciipixel = 8'hff;
				8'd08:asciipixel = 8'hff;
				8'd09:asciipixel = 8'hff;
				8'd10:asciipixel = 8'hff;
				8'd11:asciipixel = 8'h66;
				8'd12:asciipixel = 8'h66;
				8'd13:asciipixel = 8'hff;
				8'd14:asciipixel = 8'hff;
				8'd15:asciipixel = 8'hff;
				8'd16:asciipixel = 8'hff;
				8'd17:asciipixel = 8'hff;
				8'd18:asciipixel = 8'hff;
				8'd19:asciipixel = 8'hff;
				8'd20:asciipixel = 8'hff;
				8'd21:asciipixel = 8'h66;
				8'd22:asciipixel = 8'h66;
				8'd23:asciipixel = 8'hff;
				8'd24:asciipixel = 8'hff;
				8'd25:asciipixel = 8'hff;
				8'd26:asciipixel = 8'hff;
				8'd27:asciipixel = 8'hff;
				8'd28:asciipixel = 8'hff;
				8'd29:asciipixel = 8'hff;
				8'd30:asciipixel = 8'hff;
				8'd31:asciipixel = 8'h66;
				8'd32:asciipixel = 8'h66;
				8'd33:asciipixel = 8'hff;
				8'd34:asciipixel = 8'hff;
				8'd35:asciipixel = 8'hff;
				8'd36:asciipixel = 8'hff;
				8'd37:asciipixel = 8'hff;
				8'd38:asciipixel = 8'hc1;
				8'd39:asciipixel = 8'hbf;
				8'd40:asciipixel = 8'hff;
				8'd41:asciipixel = 8'h66;
				8'd42:asciipixel = 8'h66;
				8'd43:asciipixel = 8'hff;
				8'd44:asciipixel = 8'hff;
				8'd45:asciipixel = 8'hff;
				8'd46:asciipixel = 8'hd7;
				8'd47:asciipixel = 8'h4f;
				8'd48:asciipixel = 8'h1;
				8'd49:asciipixel = 8'hab;
				8'd50:asciipixel = 8'hff;
				8'd51:asciipixel = 8'h66;
				8'd52:asciipixel = 8'h66;
				8'd53:asciipixel = 8'hff;
				8'd54:asciipixel = 8'he9;
				8'd55:asciipixel = 8'h6a;
				8'd56:asciipixel = 8'h4;
				8'd57:asciipixel = 8'h3d;
				8'd58:asciipixel = 8'hc8;
				8'd59:asciipixel = 8'hff;
				8'd60:asciipixel = 8'hff;
				8'd61:asciipixel = 8'h66;
				8'd62:asciipixel = 8'h5c;
				8'd63:asciipixel = 8'h84;
				8'd64:asciipixel = 8'hd;
				8'd65:asciipixel = 8'h27;
				8'd66:asciipixel = 8'haf;
				8'd67:asciipixel = 8'hfe;
				8'd68:asciipixel = 8'hff;
				8'd69:asciipixel = 8'hff;
				8'd70:asciipixel = 8'hff;
				8'd71:asciipixel = 8'h66;
				8'd72:asciipixel = 8'h0;
				8'd73:asciipixel = 8'h16;
				8'd74:asciipixel = 8'h95;
				8'd75:asciipixel = 8'hfa;
				8'd76:asciipixel = 8'hff;
				8'd77:asciipixel = 8'hff;
				8'd78:asciipixel = 8'hff;
				8'd79:asciipixel = 8'hff;
				8'd80:asciipixel = 8'hff;
				8'd81:asciipixel = 8'h6f;
				8'd82:asciipixel = 8'h7a;
				8'd83:asciipixel = 8'hf1;
				8'd84:asciipixel = 8'hff;
				8'd85:asciipixel = 8'hff;
				8'd86:asciipixel = 8'hff;
				8'd87:asciipixel = 8'hff;
				8'd88:asciipixel = 8'hff;
				8'd89:asciipixel = 8'hff;
				8'd90:asciipixel = 8'hff;
				8'd91:asciipixel = 8'hfb;
				8'd92:asciipixel = 8'hff;
				8'd93:asciipixel = 8'hff;
				8'd94:asciipixel = 8'hff;
				8'd95:asciipixel = 8'hff;
				8'd96:asciipixel = 8'hff;
				8'd97:asciipixel = 8'hff;
				8'd98:asciipixel = 8'hff;
				8'd99:asciipixel = 8'hff;
				default:asciipixel = 0;
			endcase
		end
		else if (num == 'd11) begin // +
			case(addr)
				8'd00:asciipixel = 8'hff;
				8'd01:asciipixel = 8'hff;
				8'd02:asciipixel = 8'hff;
				8'd03:asciipixel = 8'hff;
				8'd04:asciipixel = 8'hff;
				8'd05:asciipixel = 8'hff;
				8'd06:asciipixel = 8'hff;
				8'd07:asciipixel = 8'hff;
				8'd08:asciipixel = 8'hff;
				8'd09:asciipixel = 8'hff;
				8'd10:asciipixel = 8'hff;
				8'd11:asciipixel = 8'hff;
				8'd12:asciipixel = 8'hff;
				8'd13:asciipixel = 8'hff;
				8'd14:asciipixel = 8'hcc;
				8'd15:asciipixel = 8'h0;
				8'd16:asciipixel = 8'hff;
				8'd17:asciipixel = 8'hff;
				8'd18:asciipixel = 8'hff;
				8'd19:asciipixel = 8'hff;
				8'd20:asciipixel = 8'hff;
				8'd21:asciipixel = 8'hff;
				8'd22:asciipixel = 8'hff;
				8'd23:asciipixel = 8'hff;
				8'd24:asciipixel = 8'hcc;
				8'd25:asciipixel = 8'h0;
				8'd26:asciipixel = 8'hff;
				8'd27:asciipixel = 8'hff;
				8'd28:asciipixel = 8'hff;
				8'd29:asciipixel = 8'hff;
				8'd30:asciipixel = 8'hff;
				8'd31:asciipixel = 8'hff;
				8'd32:asciipixel = 8'hff;
				8'd33:asciipixel = 8'hff;
				8'd34:asciipixel = 8'hcc;
				8'd35:asciipixel = 8'h0;
				8'd36:asciipixel = 8'hff;
				8'd37:asciipixel = 8'hff;
				8'd38:asciipixel = 8'hff;
				8'd39:asciipixel = 8'hff;
				8'd40:asciipixel = 8'hff;
				8'd41:asciipixel = 8'ha3;
				8'd42:asciipixel = 8'h66;
				8'd43:asciipixel = 8'h66;
				8'd44:asciipixel = 8'h51;
				8'd45:asciipixel = 8'h0;
				8'd46:asciipixel = 8'h66;
				8'd47:asciipixel = 8'h66;
				8'd48:asciipixel = 8'h66;
				8'd49:asciipixel = 8'hc1;
				8'd50:asciipixel = 8'hff;
				8'd51:asciipixel = 8'ha3;
				8'd52:asciipixel = 8'h66;
				8'd53:asciipixel = 8'h66;
				8'd54:asciipixel = 8'h51;
				8'd55:asciipixel = 8'h0;
				8'd56:asciipixel = 8'h66;
				8'd57:asciipixel = 8'h66;
				8'd58:asciipixel = 8'h66;
				8'd59:asciipixel = 8'hc1;
				8'd60:asciipixel = 8'hff;
				8'd61:asciipixel = 8'hff;
				8'd62:asciipixel = 8'hff;
				8'd63:asciipixel = 8'hff;
				8'd64:asciipixel = 8'hcc;
				8'd65:asciipixel = 8'h0;
				8'd66:asciipixel = 8'hff;
				8'd67:asciipixel = 8'hff;
				8'd68:asciipixel = 8'hff;
				8'd69:asciipixel = 8'hff;
				8'd70:asciipixel = 8'hff;
				8'd71:asciipixel = 8'hff;
				8'd72:asciipixel = 8'hff;
				8'd73:asciipixel = 8'hff;
				8'd74:asciipixel = 8'hcc;
				8'd75:asciipixel = 8'h0;
				8'd76:asciipixel = 8'hff;
				8'd77:asciipixel = 8'hff;
				8'd78:asciipixel = 8'hff;
				8'd79:asciipixel = 8'hff;
				8'd80:asciipixel = 8'hff;
				8'd81:asciipixel = 8'hff;
				8'd82:asciipixel = 8'hff;
				8'd83:asciipixel = 8'hff;
				8'd84:asciipixel = 8'hcc;
				8'd85:asciipixel = 8'h0;
				8'd86:asciipixel = 8'hff;
				8'd87:asciipixel = 8'hff;
				8'd88:asciipixel = 8'hff;
				8'd89:asciipixel = 8'hff;
				8'd90:asciipixel = 8'hff;
				8'd91:asciipixel = 8'hff;
				8'd92:asciipixel = 8'hff;
				8'd93:asciipixel = 8'hff;
				8'd94:asciipixel = 8'hf4;
				8'd95:asciipixel = 8'hcc;
				8'd96:asciipixel = 8'hff;
				8'd97:asciipixel = 8'hff;
				8'd98:asciipixel = 8'hff;
				8'd99:asciipixel = 8'hff;
				default:asciipixel = 0;
			endcase
		end
		else if (num == 'd14) begin // /
			case(addr)
				8'd00:asciipixel = 8'hff;
				8'd01:asciipixel = 8'hff;
				8'd02:asciipixel = 8'hff;
				8'd03:asciipixel = 8'hff;
				8'd04:asciipixel = 8'hff;
				8'd05:asciipixel = 8'hff;
				8'd06:asciipixel = 8'hff;
				8'd07:asciipixel = 8'hff;
				8'd08:asciipixel = 8'hff;
				8'd09:asciipixel = 8'hff;
				8'd10:asciipixel = 8'hff;
				8'd11:asciipixel = 8'hff;
				8'd12:asciipixel = 8'hff;
				8'd13:asciipixel = 8'hff;
				8'd14:asciipixel = 8'hff;
				8'd15:asciipixel = 8'hff;
				8'd16:asciipixel = 8'hff;
				8'd17:asciipixel = 8'hff;
				8'd18:asciipixel = 8'hff;
				8'd19:asciipixel = 8'hff;
				8'd20:asciipixel = 8'hff;
				8'd21:asciipixel = 8'hff;
				8'd22:asciipixel = 8'hff;
				8'd23:asciipixel = 8'hff;
				8'd24:asciipixel = 8'hff;
				8'd25:asciipixel = 8'hff;
				8'd26:asciipixel = 8'hff;
				8'd27:asciipixel = 8'hfb;
				8'd28:asciipixel = 8'h9a;
				8'd29:asciipixel = 8'haf;
				8'd30:asciipixel = 8'hff;
				8'd31:asciipixel = 8'hff;
				8'd32:asciipixel = 8'hff;
				8'd33:asciipixel = 8'hff;
				8'd34:asciipixel = 8'hff;
				8'd35:asciipixel = 8'hfe;
				8'd36:asciipixel = 8'hb4;
				8'd37:asciipixel = 8'h2b;
				8'd38:asciipixel = 8'hb;
				8'd39:asciipixel = 8'hbb;
				8'd40:asciipixel = 8'hff;
				8'd41:asciipixel = 8'hff;
				8'd42:asciipixel = 8'hff;
				8'd43:asciipixel = 8'hff;
				8'd44:asciipixel = 8'hcd;
				8'd45:asciipixel = 8'h42;
				8'd46:asciipixel = 8'h3;
				8'd47:asciipixel = 8'h64;
				8'd48:asciipixel = 8'he6;
				8'd49:asciipixel = 8'hff;
				8'd50:asciipixel = 8'hff;
				8'd51:asciipixel = 8'hff;
				8'd52:asciipixel = 8'he1;
				8'd53:asciipixel = 8'h5d;
				8'd54:asciipixel = 8'h1;
				8'd55:asciipixel = 8'h4a;
				8'd56:asciipixel = 8'hd4;
				8'd57:asciipixel = 8'hff;
				8'd58:asciipixel = 8'hff;
				8'd59:asciipixel = 8'hff;
				8'd60:asciipixel = 8'hff;
				8'd61:asciipixel = 8'h9c;
				8'd62:asciipixel = 8'h8;
				8'd63:asciipixel = 8'h32;
				8'd64:asciipixel = 8'hbd;
				8'd65:asciipixel = 8'hff;
				8'd66:asciipixel = 8'hff;
				8'd67:asciipixel = 8'hff;
				8'd68:asciipixel = 8'hff;
				8'd69:asciipixel = 8'hff;
				8'd70:asciipixel = 8'hff;
				8'd71:asciipixel = 8'h84;
				8'd72:asciipixel = 8'ha2;
				8'd73:asciipixel = 8'hfd;
				8'd74:asciipixel = 8'hff;
				8'd75:asciipixel = 8'hff;
				8'd76:asciipixel = 8'hff;
				8'd77:asciipixel = 8'hff;
				8'd78:asciipixel = 8'hff;
				8'd79:asciipixel = 8'hff;
				8'd80:asciipixel = 8'hff;
				8'd81:asciipixel = 8'hff;
				8'd82:asciipixel = 8'hff;
				8'd83:asciipixel = 8'hff;
				8'd84:asciipixel = 8'hff;
				8'd85:asciipixel = 8'hff;
				8'd86:asciipixel = 8'hff;
				8'd87:asciipixel = 8'hff;
				8'd88:asciipixel = 8'hff;
				8'd89:asciipixel = 8'hff;
				8'd90:asciipixel = 8'hff;
				8'd91:asciipixel = 8'hff;
				8'd92:asciipixel = 8'hff;
				8'd93:asciipixel = 8'hff;
				8'd94:asciipixel = 8'hff;
				8'd95:asciipixel = 8'hff;
				8'd96:asciipixel = 8'hff;
				8'd97:asciipixel = 8'hff;
				8'd98:asciipixel = 8'hff;
				8'd99:asciipixel = 8'hff;
				default:asciipixel = 0;
			endcase
		end
		else if (num == 'd12) begin // -
			case(addr)
				8'd00:asciipixel = 8'hff;
				8'd01:asciipixel = 8'hff;
				8'd02:asciipixel = 8'hff;
				8'd03:asciipixel = 8'hff;
				8'd04:asciipixel = 8'hff;
				8'd05:asciipixel = 8'hff;
				8'd06:asciipixel = 8'hff;
				8'd07:asciipixel = 8'hff;
				8'd08:asciipixel = 8'hff;
				8'd09:asciipixel = 8'hff;
				8'd10:asciipixel = 8'hff;
				8'd11:asciipixel = 8'hff;
				8'd12:asciipixel = 8'hff;
				8'd13:asciipixel = 8'hff;
				8'd14:asciipixel = 8'hcc;
				8'd15:asciipixel = 8'h0;
				8'd16:asciipixel = 8'hff;
				8'd17:asciipixel = 8'hff;
				8'd18:asciipixel = 8'hff;
				8'd19:asciipixel = 8'hff;
				8'd20:asciipixel = 8'hff;
				8'd21:asciipixel = 8'hff;
				8'd22:asciipixel = 8'hff;
				8'd23:asciipixel = 8'hff;
				8'd24:asciipixel = 8'hcc;
				8'd25:asciipixel = 8'h0;
				8'd26:asciipixel = 8'hff;
				8'd27:asciipixel = 8'hff;
				8'd28:asciipixel = 8'hff;
				8'd29:asciipixel = 8'hff;
				8'd30:asciipixel = 8'hff;
				8'd31:asciipixel = 8'hff;
				8'd32:asciipixel = 8'hff;
				8'd33:asciipixel = 8'hff;
				8'd34:asciipixel = 8'hcc;
				8'd35:asciipixel = 8'h0;
				8'd36:asciipixel = 8'hff;
				8'd37:asciipixel = 8'hff;
				8'd38:asciipixel = 8'hff;
				8'd39:asciipixel = 8'hff;
				8'd40:asciipixel = 8'hff;
				8'd41:asciipixel = 8'hff;
				8'd42:asciipixel = 8'hff;
				8'd43:asciipixel = 8'hff;
				8'd44:asciipixel = 8'hcc;
				8'd45:asciipixel = 8'h0;
				8'd46:asciipixel = 8'hff;
				8'd47:asciipixel = 8'hff;
				8'd48:asciipixel = 8'hff;
				8'd49:asciipixel = 8'hff;
				8'd50:asciipixel = 8'hff;
				8'd51:asciipixel = 8'hff;
				8'd52:asciipixel = 8'hff;
				8'd53:asciipixel = 8'hff;
				8'd54:asciipixel = 8'hcc;
				8'd55:asciipixel = 8'h0;
				8'd56:asciipixel = 8'hff;
				8'd57:asciipixel = 8'hff;
				8'd58:asciipixel = 8'hff;
				8'd59:asciipixel = 8'hff;
				8'd60:asciipixel = 8'hff;
				8'd61:asciipixel = 8'hff;
				8'd62:asciipixel = 8'hff;
				8'd63:asciipixel = 8'hff;
				8'd64:asciipixel = 8'hcc;
				8'd65:asciipixel = 8'h0;
				8'd66:asciipixel = 8'hff;
				8'd67:asciipixel = 8'hff;
				8'd68:asciipixel = 8'hff;
				8'd69:asciipixel = 8'hff;
				8'd70:asciipixel = 8'hff;
				8'd71:asciipixel = 8'hff;
				8'd72:asciipixel = 8'hff;
				8'd73:asciipixel = 8'hff;
				8'd74:asciipixel = 8'hcc;
				8'd75:asciipixel = 8'h0;
				8'd76:asciipixel = 8'hff;
				8'd77:asciipixel = 8'hff;
				8'd78:asciipixel = 8'hff;
				8'd79:asciipixel = 8'hff;
				8'd80:asciipixel = 8'hff;
				8'd81:asciipixel = 8'hff;
				8'd82:asciipixel = 8'hff;
				8'd83:asciipixel = 8'hff;
				8'd84:asciipixel = 8'hcc;
				8'd85:asciipixel = 8'h0;
				8'd86:asciipixel = 8'hff;
				8'd87:asciipixel = 8'hff;
				8'd88:asciipixel = 8'hff;
				8'd89:asciipixel = 8'hff;
				8'd90:asciipixel = 8'hff;
				8'd91:asciipixel = 8'hff;
				8'd92:asciipixel = 8'hff;
				8'd93:asciipixel = 8'hff;
				8'd94:asciipixel = 8'hf4;
				8'd95:asciipixel = 8'hcc;
				8'd96:asciipixel = 8'hff;
				8'd97:asciipixel = 8'hff;
				8'd98:asciipixel = 8'hff;
				8'd99:asciipixel = 8'hff;
				default:asciipixel = 0;
			endcase
		end
        else begin
            asciipixel = 8'd0;
        end
endmodule