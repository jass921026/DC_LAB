`timescale 1ns/1ns

module wt_mem7 #(parameter ADDR_WIDTH = 11, DATA_WIDTH = 144, DEPTH = 76) (
input wire clk,
input wire [ADDR_WIDTH-1:0] addr_a, 
input wire [ADDR_WIDTH-1:0] addr_b, 
output reg [DATA_WIDTH-1:0] q_a,
output reg [DATA_WIDTH-1:0] q_b
);

reg [DATA_WIDTH-1:0] mem [0:DEPTH-1];

initial begin
mem[0] = 144'h118b15aa0368f8e81ad60baeff320bb3f4fc;
mem[1] = 144'hee93ef0ef705fbda0122fea50f7bf69cf8fa;
mem[2] = 144'hf7d5f8b0f8cafc32fe9601dffe55fa7cffa0;
mem[3] = 144'hfd3c04a0fd1403940526fbab013104a5fe74;
mem[4] = 144'hf936002dfffefbd006e3febaff29fc9cfcc2;
mem[5] = 144'h016903dffd01ff6ffbd5fdf9fe97ffcb052e;
mem[6] = 144'hfe22f793f5e2021304f4fec6fe600061fbce;
mem[7] = 144'h0090033a0532012b00c4fcb4fb88fdbbfb18;
mem[8] = 144'hfab9fe600115fd75fc9dfeb8050501310058;
mem[9] = 144'h0323fb9f004202bafb7cfc8e044e02610402;
mem[10] = 144'hfcadfac7fb22f91cfd6f014ffb7afd330507;
mem[11] = 144'hff85fe87031afe7bfaef003d03910254fce8;
mem[12] = 144'h027eff44ffc1032afd00fe4705d605cb024f;
mem[13] = 144'hfd57fe09fd4eff95fc25fad0fe720235039b;
mem[14] = 144'hf7b7f997f644fc880205fa02052a05acfda0;
mem[15] = 144'h054dfb74fcd702240126fe10fc37fee8fd63;
mem[16] = 144'hf7abfa4f074af2bbffd90602feb8040602b3;
mem[17] = 144'h03c40111fec4fb75febe012afc9a000dfbc5;
mem[18] = 144'hfc5ffa3afb07fc61fe90fe430387ff5e032a;
mem[19] = 144'hfcc90154fe51049202f8fc00004a028a02bf;
mem[20] = 144'hf71cfef2f5e2ffc8fbd8f75f017d005b01b9;
mem[21] = 144'h017900d7ffca01eafe08fc50fef6024cfc1e;
mem[22] = 144'h04b3fec2fbb000d305abfde607df0521ff2e;
mem[23] = 144'h00b40364fb0affa9043bfecf031dfefa047f;
mem[24] = 144'hff80f973f924012ffdf1007900450281fba9;
mem[25] = 144'h011cff30fd4dfb13fe9afd0efd1cfb970029;
mem[26] = 144'hff86f8e5fbf3fec6013c03e70149003d0822;
mem[27] = 144'hfc46fd670131febafc1efe60fe38fc91ffec;
mem[28] = 144'hf5d4f64cffe9fe71fa5ffebbfb6b05f20101;
mem[29] = 144'h02ab040bfab8ffa5fc86038a004d041bffb2;
mem[30] = 144'h0518fdc9009206bd00e2fed500dc038906a4;
mem[31] = 144'hfc340271fee9fe2102f5fceaff7604fefac0;
mem[32] = 144'hfbe000360079fb120081fa11039a0432f98b;
mem[33] = 144'h04adfca1fde3051104f1fdc4fc7d04b1fe09;
mem[34] = 144'hfde0f5affb6bfca3028d02f8fffffe65fc3d;
mem[35] = 144'h00d9010704c4fdfe0364feb5045afe4f053b;
mem[36] = 144'h0272fc6ef975fc3df8fb012fffe3fdd6ffd0;
mem[37] = 144'hffe2045e022c0472fb26fcc4fb66ff780064;
mem[38] = 144'hf834fe18f5090192036cf8f4fe17035efbb6;
mem[39] = 144'hff9ffe620338fdf6fb1a047cfe1c00dcfb46;
mem[40] = 144'hf9f3f891f6b7ff7dfbcbff48fdc9033902ed;
mem[41] = 144'h02e1fbabfd27fd720468fecdfb7601dffae1;
mem[42] = 144'hfcbdfd8df419fb97000401d0fe9902a6faca;
mem[43] = 144'h055501e7fd55ffb104e4fb35016efc15fbde;
mem[44] = 144'h0925038603850232fe72ff5f017d06c603d0;
mem[45] = 144'hfce9fecc001cff08013200d50388028b0306;
mem[46] = 144'h05f1020b09d90381feae043dff8501d50607;
mem[47] = 144'hfb43fc23fb3efc8a010d02f80093017aff10;
mem[48] = 144'h0713fefe01b90048022dfbf706f5064d021e;
mem[49] = 144'hfbd3fd180126fffeff5803950068ffcc0543;
mem[50] = 144'hfe8a01c902effa5bfd3303dcfcbcfc08fa56;
mem[51] = 144'hff1402790130fcdc03ef0295031604b20383;
mem[52] = 144'hffc5ff56052100300447ff3efe47fc8a06fd;
mem[53] = 144'h004afcccfbf6016e04b1fdb4fd06ffba04ea;
mem[54] = 144'hfbd9fe58fdc7fdab03a4fee1fc0f01f30203;
mem[55] = 144'h0029fd15fc3aff31001efb66fc6eff03ff73;
mem[56] = 144'h0ada0bb10ac5039b09c206a4ff84fd040246;
mem[57] = 144'h0003fbf204a6ff08028b00d4049400500335;
mem[58] = 144'h006604e1035506dd048105d2fcf601a8fc63;
mem[59] = 144'h02d8fcfc040a046e02dd0175fff9fbd6fdd1;
mem[60] = 144'hfe04ff8cfab5f7abfb0cfaeafe2b06affd5b;
mem[61] = 144'hfc98ffc3fcbcfee302bcfbc3ffb0fd53ff0d;
mem[62] = 144'hfee0fcf7fcb0f7d2ff88ffe5fec90242022f;
mem[63] = 144'hfd91fdb5fec7fc2b005d04d2ff69015e0361;
mem[64] = 144'hf3b8f673f4c4f8700007fe010117016c03eb;
mem[65] = 144'h0434019103d8fe6d029802a0ffd302aefbdb;
mem[66] = {16'hfce4, 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000};
mem[67] = {16'hf73f, 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000};
mem[68] = {16'hfdd5, 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000};
mem[69] = {16'hfcf0, 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000};
mem[70] = {16'hfd58, 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000};
mem[71] = {16'h0b3d, 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000};
mem[72] = {16'hf830, 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000};
mem[73] = {16'h0597, 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000};
mem[74] = {16'hf8bc, 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000};
mem[75] = {16'h0927, 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000};
end

always @ (posedge clk) begin
	q_a <= mem[addr_a];
end

always @ (posedge clk) begin
	q_b <= mem[addr_b];
end

endmodule