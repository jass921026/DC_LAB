module CNN_test
#(
    parameter GS_BITS = 8, 
    parameter BCD_BITS = 4 
)
(
    input clk,
    input rst,
    output reg [GS_BITS-1:0] pixel_i,
    output reg pixel_i_valid
);
    logic [19:0] count_time;
    logic [4:0] digit;
    logic [4:0] x, y;

    //counter
    Counter #(
        .WIDTH(20),
        .MAX_COUNT(500000)
    ) counter (
        .clk(clk),
        .rst_n(rst),
        .enable(1'b1),
        .count(count_time)
    );

    //digit
    Counter #(
        .WIDTH(4),
        .MAX_COUNT(9)
    ) digit_counter (
        .clk(clk),
        .rst_n(rst),
        .enable(count_time == 20'd499999),
        .count(digit)
    );

    //xy  
    Counter #(
        .WIDTH(5),
        .MAX_COUNT(29)
    ) x_counter (
        .clk(clk),
        .rst_n(count_time == 20'd499999),
        .enable(1'b1),
        .count(x)
    );
    Counter #(
        .WIDTH(5),
        .MAX_COUNT(29)
    ) y_counter (
        .clk(clk),
        .rst_n(count_time == 20'd499999),
        .enable(x == 29),
        .count(y)
    );

    //pixel

    logic [29:0][29:0] digit_1 = '{
            30'b000000000000000000000000000000,
            30'b000000000000000000000000000000,
            30'b000000000000000000000000000000,
            30'b000000000000000000000000000000,
            30'b000000000000011000000000000000,
            30'b000000011111111000000000000000,
            30'b000000000000011000000000000000,
            30'b000000000000011000000000000000,
            30'b000000000000011000000000000000,
            30'b000000000000011000000000000000,
            30'b000000000000011000000000000000,
            30'b000000000000011000000000000000,
            30'b000000000000011000000000000000,
            30'b000000000000011000000000000000,
            30'b000000000000011000000000000000,
            30'b000000000000011000000000000000,
            30'b000000000000011000000000000000,
            30'b000000000000011000000000000000,
            30'b000000000000011000000000000000,
            30'b000000000000011000000000000000,
            30'b000000000000011000000000000000,
            30'b000000000000011000000000000000,
            30'b000000111111111111111110000000,
            30'b000000000000000000000000000000,
            30'b000000000000000000000000000000,
            30'b000000000000000000000000000000,
            30'b000000000000000000000000000000,
            30'b000000000000000000000000000000,
            30'b000000000000000000000000000000,
            30'b000000000000000000000000000000
    };

    assign pixel_i = digit_1[x][y] ? 8'b11111111 : 8'b00000000;
    assign pixel_i_valid = count_time < 20'd900 ? 1 : 0;


endmodule