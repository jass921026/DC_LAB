module Magic_mask
(
    input [3:0] idx,
    output [29:0][29:0] mask 
);

    logic [29:0][29:0] digit_blank = '{
            30'b000000000000000000000000000000,
            30'b000000000000000000000000000000,
            30'b000000000000000000000000000000,
            30'b000000000000000000000000000000,
            30'b000000000000000000000000000000,
            30'b000000000000000000000000000000,
            30'b000000000000000000000000000000,
            30'b000000000000000000000000000000,
            30'b000000000000000000000000000000,
            30'b000000000000000000000000000000,
            30'b000000000000000000000000000000,
            30'b000000000000000000000000000000,
            30'b000000000000000000000000000000,
            30'b000000000000000000000000000000,
            30'b000000000000000000000000000000,
            30'b000000000000000000000000000000,
            30'b000000000000000000000000000000,
            30'b000000000000000000000000000000,
            30'b000000000000000000000000000000,
            30'b000000000000000000000000000000,
            30'b000000000000000000000000000000,
            30'b000000000000000000000000000000,
            30'b000000000000000000000000000000,
            30'b000000000000000000000000000000,
            30'b000000000000000000000000000000,
            30'b000000000000000000000000000000,
            30'b000000000000000000000000000000,
            30'b000000000000000000000000000000,
            30'b000000000000000000000000000000,
            30'b000000000000000000000000000000
    };
    
    logic [29:0][29:0] digit_0 = '{
            30'b000000000000000000000000000000,
            30'b000000000000000000000000000000,
            30'b000000000000000000000000000000,
            30'b000000000000000000000000000000,
            30'b000000000000000000000000000000,
            30'b000000000000000000000000000000,
            30'b000000000000000000000000000000,
            30'b000000000000000000000000000000,
            30'b000000000000000000000000000000,
            30'b000000000000000000000000000000,
            30'b000000000000000000000000000000,
            30'b000000000000000000000000000000,
            30'b000000000000000000000000000000,
            30'b000000000000000000000000000000,
            30'b000000000000000000000000000000,
            30'b000000000000000000000000000000,
            30'b000000000000000000000000000000,
            30'b000000000000000000000000000000,
            30'b000000000000000000000000000000,
            30'b000000000000000000000000000000,
            30'b000000000000000000000000000000,
            30'b000000000000000000000000000000,
            30'b000000000000000000000000000000,
            30'b000000000000000000000000000000,
            30'b000000000000000000000000000000,
            30'b000000000000000000000000000000,
            30'b000000000000000000000000000000,
            30'b000000000000000000000000000000,
            30'b000000000000000000000000000000,
            30'b000000000000000000000000000000
    };

    logic [29:0][29:0] digit_1 = '{
            30'b000000000000000000000000000000,
            30'b000000000000000000000000000000,
            30'b000000000000000000000000000000,
            30'b000000000000000000000000000000,
            30'b000000000000000000000000000000,
            30'b000000000000000000000000000000,
            30'b000000000000000000000000000000,
            30'b000000000000000000000000000000,
            30'b000000000000000000000000000000,
            30'b000000000000000000000000000000,
            30'b000000000000000000000000000000,
            30'b000000000000000000000000000000,
            30'b000000000000000000000000000000,
            30'b000000000000000000000000000000,
            30'b000000000000000000000000000000,
            30'b000000000000000000000000000000,
            30'b000000000000000000000000000000,
            30'b000000000000000000000000000000,
            30'b000000000000000000000000000000,
            30'b000000000000000000000000000000,
            30'b000000000000000000000000000000,
            30'b000000000000000000000000000000,
            30'b000000000000000000000000000000,
            30'b000000000000000000000000000000,
            30'b000000000000000000000000000000,
            30'b000000000000000000000000000000,
            30'b000000000000000000000000000000,
            30'b000000000000000000000000000000,
            30'b000000000000000000000000000000,
            30'b000000000000000000000000000000
    };

    logic [29:0][29:0] digit_2 = '{
            30'b000000000000000000000000000000,
            30'b000000000000000000000000000000,
            30'b000000000000000000000000000000,
            30'b000000000000000000000000000000,
            30'b000000000000000000000000000000,
            30'b000000000000000000000000000000,
            30'b000000000000000000000000000000,
            30'b000000000000000000000000000000,
            30'b000000000000000000000000000000,
            30'b000000000000000000000000000000,
            30'b000000000000000000000000000000,
            30'b000000000000000000000000000000,
            30'b000000000000000000000000000000,
            30'b000000000000000000000000000000,
            30'b000000000000000000000000000000,
            30'b000000000000000000000000000000,
            30'b000000000000000000000000000000,
            30'b000000000000000000000000000000,
            30'b000000000000000000000000000000,
            30'b000000000000000000000000000000,
            30'b000000000000000000000000000000,
            30'b000000000000000000000000000000,
            30'b000000000000000000000000000000,
            30'b000000000000000000000000000000,
            30'b000000000000000000000000000000,
            30'b000000000000000000000000000000,
            30'b000000000000000000000000000000,
            30'b000000000000000000000000000000,
            30'b000000000000000000000000000000,
            30'b000000000000000000000000000000
    };

    logic [29:0][29:0] digit_3 = '{
            30'b000000000000000000000000000000,
            30'b000000000000000000000000000000,
            30'b000000000000000000000000000000,
            30'b000000000000000000000000000000,
            30'b000000000000000000000000000000,
            30'b000000000000000000000000000000,
            30'b000000000000000000000000000000,
            30'b000000000000000000000000000000,
            30'b000000000000000000000000000000,
            30'b000000000000000000000000000000,
            30'b000000000000000000000000000000,
            30'b000000000000000000000000000000,
            30'b000000000000000000000000000000,
            30'b000000000000000000000000000000,
            30'b000000000000000000000000000000,
            30'b000000000000000000000000000000,
            30'b000000000000000000000000000000,
            30'b000000000000000000000000000000,
            30'b000000000000000000000000000000,
            30'b000000000000000000000000000000,
            30'b000000000000000000000000000000,
            30'b000000000000000000000000000000,
            30'b000000000000000000000000000000,
            30'b000000000000000000000000000000,
            30'b000000000000000000000000000000,
            30'b000000000000000000000000000000,
            30'b000000000000000000000000000000,
            30'b000000000000000000000000000000,
            30'b000000000000000000000000000000,
            30'b000000000000000000000000000000
    };

    logic [29:0][29:0] digit_4 = '{
            30'b000000000000000000000000000000,
            30'b000000000000000000000000000000,
            30'b000000000000000000000000000000,
            30'b000000000000000000000000000000,
            30'b000000000000000000000000000000,
            30'b000000000000000000000000000000,
            30'b000000000000000000000000000000,
            30'b000000000000000000000000000000,
            30'b000000000000000000000000000000,
            30'b000000000000000000000000000000,
            30'b000000000000000000000000000000,
            30'b000000000000000000000000000000,
            30'b000000000000000000000000000000,
            30'b000000000000000000000000000000,
            30'b000000000000000000000000000000,
            30'b000000000000000000000000000000,
            30'b000000000000000000000000000000,
            30'b000000000000000000000000000000,
            30'b000000000000000000000000000000,
            30'b000000000000000000000000000000,
            30'b000000000000000000000000000000,
            30'b000000000000000000000000000000,
            30'b000000000000000000000000000000,
            30'b000000000000000000000000000000,
            30'b000000000000000000000000000000,
            30'b000000000000000000000000000000,
            30'b000000000000000000000000000000,
            30'b000000000000000000000000000000,
            30'b000000000000000000000000000000,
            30'b000000000000000000000000000000
    };

    logic [29:0][29:0] digit_5 = '{
            30'b000000000000000000000000000000,
            30'b000000000000000000000000000000,
            30'b000000000000000000000000000000,
            30'b000000000000000000000000000000,
            30'b000000000000000000000000000000,
            30'b000000000000000000000000000000,
            30'b000000000000000000000000000000,
            30'b000000000000000000000000000000,
            30'b000000000000000000000000000000,
            30'b000000000000000000000000000000,
            30'b000000000000000000000000000000,
            30'b000000000000000000000000000000,
            30'b000000000000000000000000000000,
            30'b000000000000000000000000000000,
            30'b000000000000000000000000000000,
            30'b000000000000000000000000000000,
            30'b000000000000000000000000000000,
            30'b000000000000000000000000000000,
            30'b000000000000000000000000000000,
            30'b000000000000000000000000000000,
            30'b000000000000000000000000000000,
            30'b000000000000000000000000000000,
            30'b000000000000000000000000000000,
            30'b000000000000000000000000000000,
            30'b000000000000000000000000000000,
            30'b000000000000000000000000000000,
            30'b000000000000000000000000000000,
            30'b000000000000000000000000000000,
            30'b000000000000000000000000000000,
            30'b000000000000000000000000000000
    };

    logic [29:0][29:0] digit_6 = '{
            30'b000000000000000000000000000000,
            30'b000000000000000000000000000000,
            30'b000000000000000000000000000000,
            30'b000000000000000000000000000000,
            30'b000000000000000000000000000000,
            30'b000000000000000000000000000000,
            30'b000000000000000000000000000000,
            30'b000000000000000000000000000000,
            30'b000000000000000000000000000000,
            30'b000000000000000000000000000000,
            30'b000000000000000000000000000000,
            30'b000000000000000000000000000000,
            30'b000000000000000000000000000000,
            30'b000000000000000000000000000000,
            30'b000000000000000000000000000000,
            30'b000000000000000000000000000000,
            30'b000000000000000000000000000000,
            30'b000000000000000000000000000000,
            30'b000000000000000000000000000000,
            30'b000000000000000000000000000000,
            30'b000000000000000000000000000000,
            30'b000000000000000000000000000000,
            30'b000000000000000000000000000000,
            30'b000000000000000000000000000000,
            30'b000000000000000000000000000000,
            30'b000000000000000000000000000000,
            30'b000000000000000000000000000000,
            30'b000000000000000000000000000000,
            30'b000000000000000000000000000000,
            30'b000000000000000000000000000000
    };

    logic [29:0][29:0] digit_7 = '{
            30'b000000000000000000000000000000,
            30'b000000000000000000000000000000,
            30'b000000000000000000000000000000,
            30'b000000000000000000000000000000,
            30'b000000000000000000000000000000,
            30'b000000000000000000000000000000,
            30'b000000000000000000000000000000,
            30'b000000000000000000000000000000,
            30'b000000000000000000000000000000,
            30'b000000000000000000000000000000,
            30'b000000000000000000000000000000,
            30'b000000000000000000000000000000,
            30'b000000000000000000000000000000,
            30'b000000000000000000000000000000,
            30'b000000000000000000000000000000,
            30'b000000000000000000000000000000,
            30'b000000000000000000000000000000,
            30'b000000000000000000000000000000,
            30'b000000000000000000000000000000,
            30'b000000000000000000000000000000,
            30'b000000000000000000000000000000,
            30'b000000000000000000000000000000,
            30'b000000000000000000000000000000,
            30'b000000000000000000000000000000,
            30'b000000000000000000000000000000,
            30'b000000000000000000000000000000,
            30'b000000000000000000000000000000,
            30'b000000000000000000000000000000,
            30'b000000000000000000000000000000,
            30'b000000000000000000000000000000
    };

    logic [29:0][29:0] digit_8 = '{
            30'b000000000000000000000000000000,
            30'b000000000000000000000000000000,
            30'b000000000000000000000000000000,
            30'b000000000000000000000000000000,
            30'b000000000000000000000000000000,
            30'b000000000000000000000000000000,
            30'b000000000000000000000000000000,
            30'b000000000000000000000000000000,
            30'b000000000000000000000000000000,
            30'b000000000000000000000000000000,
            30'b000000000000000000000000000000,
            30'b000000000000000000000000000000,
            30'b000000000000000000000000000000,
            30'b000000000000000000000000000000,
            30'b000000000000000000000000000000,
            30'b000000000000000000000000000000,
            30'b000000000000000000000000000000,
            30'b000000000000000000000000000000,
            30'b000000000000000000000000000000,
            30'b000000000000000000000000000000,
            30'b000000000000000000000000000000,
            30'b000000000000000000000000000000,
            30'b000000000000000000000000000000,
            30'b000000000000000000000000000000,
            30'b000000000000000000000000000000,
            30'b000000000000000000000000000000,
            30'b000000000000000000000000000000,
            30'b000000000000000000000000000000,
            30'b000000000000000000000000000000,
            30'b000000000000000000000000000000
    };

    logic [29:0][29:0] digit_9 = '{
            30'b000000000000000000000000000000,
            30'b000000000000000000000000000000,
            30'b000000000000000000000000000000,
            30'b000000000000000000000000000000,
            30'b000000000000000000000000000000,
            30'b000000000000000000000000000000,
            30'b000000000000000000000000000000,
            30'b000000000000000000000000000000,
            30'b000000000000000000000000000000,
            30'b000000000000000000000000000000,
            30'b000000000000000000000000000000,
            30'b000000000000000000000000000000,
            30'b000000000000000000000000000000,
            30'b000000000000000000000000000000,
            30'b000000000000000000000000000000,
            30'b000000000000000000000000000000,
            30'b000000000000000000000000000000,
            30'b000000000000000000000000000000,
            30'b000000000000000000000000000000,
            30'b000000000000000000000000000000,
            30'b000000000000000000000000000000,
            30'b000000000000000000000000000000,
            30'b000000000000000000000000000000,
            30'b000000000000000000000000000000,
            30'b000000000000000000000000000000,
            30'b000000000000000000000000000000,
            30'b000000000000000000000000000000,
            30'b000000000000000000000000000000,
            30'b000000000000000000000000000000,
            30'b000000000000000000000000000000
    };

    always_comb begin
        case (idx)
            4'd0: mask = digit_0;
            4'd1: mask = digit_1;
            4'd2: mask = digit_2;
            4'd3: mask = digit_3;
            4'd4: mask = digit_4;
            4'd5: mask = digit_5;
            4'd6: mask = digit_6;
            4'd7: mask = digit_7;
            4'd8: mask = digit_8;
            4'd9: mask = digit_9;
            default: mask = digit_blank;
        endcase
    end

endmodule