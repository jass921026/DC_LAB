`timescale 1ns/1ns

module wt_mem5 #(parameter ADDR_WIDTH = 11, DATA_WIDTH = 144, DEPTH = 76) (
input wire clk,
input wire [ADDR_WIDTH-1:0] addr_a, 
input wire [ADDR_WIDTH-1:0] addr_b, 
output reg [DATA_WIDTH-1:0] q_a,
output reg [DATA_WIDTH-1:0] q_b
);

reg [DATA_WIDTH-1:0] mem [0:DEPTH-1];

initial begin
mem[0] = 144'hf5b009cffbc00693108ff3d511170c9d1f70;
mem[1] = 144'h127818b205f20a8c123b1b330388ff6df62d;
mem[2] = 144'hfe790641fb7cfaca02cd03e6f7a0fc65fb4c;
mem[3] = 144'hfcd0010df8a40cbe05160422002e07a00223;
mem[4] = 144'h0480ff9f017afb24feb500a8f82afc8cf6a2;
mem[5] = 144'h080405e5fe2801d80b3c0851023efef602b9;
mem[6] = 144'h0526fd2d04980367fae4fd65fab9fb67f6d4;
mem[7] = 144'h05cb047901350aba0b5f073800090922040a;
mem[8] = 144'h009603d600c60680028f00aafe3b0246037a;
mem[9] = 144'hf43df1b8f25bf4e3f9e2fc1f0ae00a91068b;
mem[10] = 144'hf798f9bfff2a0122fe6401eb056804e90449;
mem[11] = 144'hfa25f503ff5eec92fa1401a0f6ca00f30de6;
mem[12] = 144'hfe8d033cfda903de0029046c0a890b5c06a8;
mem[13] = 144'hf96ef6a7f2baf607f558fd3d052100a60231;
mem[14] = 144'hff0e04abfce1021d0518fc26fca6fbb8f9f1;
mem[15] = 144'hf3ebf78101eefe5e050708870abd05630141;
mem[16] = 144'hf16800620100f582fa2e00ca014efd95f712;
mem[17] = 144'hf61b027d0a61f32cfe960feaf6d6fd170a6a;
mem[18] = 144'h00eaff83fc22fd1d01d5fca20194fd74f773;
mem[19] = 144'hf742f35bfa01fe9208eb006706900844ffb1;
mem[20] = 144'hfd3bfe0cf943057b05f3ff83f63d0008fab3;
mem[21] = 144'hfb2c0083fae20aa00d6f00d1096609380634;
mem[22] = 144'h08e6064501690a3e0623024c09f900a5016a;
mem[23] = 144'h0080ff98f804ff35fa18f0360466ffd9f1dd;
mem[24] = 144'h030efdd5fe81fd36ff1dff26fdee028bfd3e;
mem[25] = 144'hfdbefc58fcdcfc9b028100080484fa5ffe50;
mem[26] = 144'hfb2702ff01cf08ca05bd062f025cff110582;
mem[27] = 144'hf38decf4f7b9f9e5fde4ff1e0d9804b40680;
mem[28] = 144'hfc51fce4011cfb7bfda1fbb5fee400b70211;
mem[29] = 144'hf3c8fdcffa14fb84fbe905c60368098f017c;
mem[30] = 144'h052bfcac071f0700019a074b0295069708cb;
mem[31] = 144'hf336f411f4b6f089f396fd24fe3cfda6086b;
mem[32] = 144'h0129024e02d6fda80261fd2afc35fa30f7b9;
mem[33] = 144'h0240faf3fa60fecf045cff4400d709900259;
mem[34] = 144'hff5cff2f04edff090122fb6cf79dfa8dfc0b;
mem[35] = 144'hf8130221f84607a2066604020227021f027b;
mem[36] = 144'hfbf2feaa013003eb05b801f306c903450934;
mem[37] = 144'hfcd7f51dfa8af8090051f9a6fe5a08210ae1;
mem[38] = 144'h065c006ffc62017005b605fbf9b1fc3bf7f3;
mem[39] = 144'hfc25ff5bf064059d05810635fe2504fc0187;
mem[40] = 144'hfee90193fe1d020e02b80237fc7b037bfef6;
mem[41] = 144'hf85cf759f862fc4bfeb105a803300c5b08ab;
mem[42] = 144'h0550048dfe11048002f60530031c02e3fee8;
mem[43] = 144'hfa21f7e7fc9803430245fca601670d4b0804;
mem[44] = 144'hffa407d40265087d0593fe560805081f055a;
mem[45] = 144'h0d9f0277fe9c0481015ff2f20575fe4bf58e;
mem[46] = 144'h0125018001dcfa8dff690b04fc2b044403fe;
mem[47] = 144'hf516fb6208ecef9ff3a809ebeedefc1e027e;
mem[48] = 144'h0488fd6dff70079701b1020d04f503f7fba8;
mem[49] = 144'h082903eaf5b90b950243f73a04c200b3f808;
mem[50] = 144'h00f8fa88fb7cf9a2ffc8faeefb5002b7fa43;
mem[51] = 144'h040201ab039c01920324ffe90169fea4fa7e;
mem[52] = 144'h0160017503fffd5a02ef0420fd92018b05f9;
mem[53] = 144'hfcb3fdd502c2f90bfa2408ddf4bffb2502e8;
mem[54] = 144'hfd4a00ed0254fee4fa7801c503cdfbd4ff2e;
mem[55] = 144'hfbc4ff4dfc35031b02defe2dfc2affc7fb99;
mem[56] = 144'h079a086a06ddf78df756f903fa5bfbb4fcc0;
mem[57] = 144'h11cd131b0f88057c09020dd4f014f18ef722;
mem[58] = 144'h03fa0752fcf7fa39fd37fe81efe8f8b8f3c4;
mem[59] = 144'h073405fe06f4085c0cab0a24ffaa0110fe56;
mem[60] = 144'hffb0fe79ff28026b05de0018fd6cfd730099;
mem[61] = 144'hfb92fe2bf8a5f749ff490481078a03e30565;
mem[62] = 144'hfd31fc8efbf4fdec04b30143fee7fae2fa27;
mem[63] = 144'hf6affce1fde807dd028302ba054704d9fec5;
mem[64] = 144'h02a8fee503b00028003cfbd9fc00fe11f845;
mem[65] = 144'hf94afd81f78701c700ed00fc01a40a7f08c0;
mem[66] = 144'hff1603e9f84e0160fa56fa48f6bf066c010f;
mem[67] = 144'h09c8ff820939fedd0619f86b05ba07ecf59c;
mem[68] = 144'h017bfcd80731092e07e3027bfb72f530fe22;
mem[69] = 144'hfdc2ff2c0646f6840612fedf09a0f818fb96;
mem[70] = 144'hfd60fe30fdc7fd5b0380051ff9da01cdf935;
mem[71] = 144'h05bf01db05d3f575044306b2ff0ffd4b06f8;
mem[72] = 144'hf7d5f840fbc5002c08100533086006b8062e;
mem[73] = 144'h028efd0308370ab2f6c2f9940869032e0815;
mem[74] = 144'h0722061b063ef6940539056ff4d4067bfc47;
mem[75] = 144'h00ea0660f546f96203c4037cffa60774f384;
end

always @ (posedge clk) begin
	q_a <= mem[addr_a];
end

always @ (posedge clk) begin
	q_b <= mem[addr_b];
end

endmodule