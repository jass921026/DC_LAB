`timescale 1ns/1ns

module wt_fc1_mem3 #(parameter ADDR_WIDTH = 11, DATA_WIDTH = 144, DEPTH = 1024) (
input wire clk,
input wire [ADDR_WIDTH-1:0] addr_a, 
input wire [ADDR_WIDTH-1:0] addr_b, 
output reg [DATA_WIDTH-1:0] q_a,
output reg [DATA_WIDTH-1:0] q_b
);

reg [DATA_WIDTH-1:0] mem [0:DEPTH-1];

initial begin
mem[0] = 144'h022d03e901f7039001de020eff44016302fb;
mem[1] = 144'h03b6009f006a02a50281014b000cfe88023c;
mem[2] = 144'hfd20ff600272021f0180fc28fb62fe0afe1a;
mem[3] = 144'h026f02cc033604fb01910035fbdaff1e00c1;
mem[4] = 144'h02af014d0014031d00b500ccfe96015800a8;
mem[5] = 144'hfb08ff01fe88fef4fcd1fe45fca3fe0ffe0c;
mem[6] = 144'h0218035c0264fdbcfff4001cfd22ff960108;
mem[7] = 144'hfcc8fe800007ff96ff3bff030016fa28fe0d;
mem[8] = 144'h0020011202de04b2013d0166fd0bff440174;
mem[9] = 144'h008c0213006f026a014cfea8fe7efe170177;
mem[10] = 144'h026e01c40172013a0041fd7afe2fffec02dc;
mem[11] = 144'hfa11f660fa7602800211fc06fb13ffe5fdde;
mem[12] = 144'hff88fdb0011f01b8ff0500a100cffeb700e3;
mem[13] = 144'h0155ffd300ac0075fee1fe240034ff83fffe;
mem[14] = 144'h009e03f80228024b047c01a301d0006e010c;
mem[15] = 144'h0021006d028202b2040cffb4ffcaff000394;
mem[16] = 144'hffabfecffeacfe96ffc9fdc40177fe5d0041;
mem[17] = 144'hfeeffe0dfff6ff06004cfdc4ff4001310163;
mem[18] = 144'hfee100d400db00d80238fe1b0012ff70fe40;
mem[19] = 144'hfded01b9ffa50106ffc300e60091ff8dffd5;
mem[20] = 144'h003c0059fee2010fffd5fefdfffd006cfff6;
mem[21] = 144'h00a80067ffb5012dffd60047fdec01680081;
mem[22] = 144'h02120138ffd200570044ff50ffa3005efe57;
mem[23] = 144'hfef4002afdfdffccfea7ff27019200260159;
mem[24] = 144'hfe7affa600cf005cfe58ff9a012fff21017d;
mem[25] = 144'hfec7017200b100effec90219fed3fee701aa;
mem[26] = 144'h01c9fe170102ffcaff38ff74fdef014aff3d;
mem[27] = 144'h013ffe85ff6a0148fe450098fec1ff15ff13;
mem[28] = 144'hff4e0077017900260161fe8e011dfe3801dc;
mem[29] = 144'h00f9ff4d01cd0173ffc5000f011f0106011e;
mem[30] = 144'hfe65007bfebb00cc00cc0090ff17fedcfef5;
mem[31] = 144'hfdd1fffaff80ff3cfe22ffd0fdc700eafe36;
mem[32] = 144'hff2eff2dff33fe32fe1cfebafe0e0049017d;
mem[33] = 144'hfde7ff55feb100ac017600e9001f011b00cc;
mem[34] = 144'h00adfe8800b7fe370109ff48006eff720163;
mem[35] = 144'h000bfee00171ff3ffe2100dcfe5500470123;
mem[36] = 144'h00ae0090ffb8fe42feae01370032001f0181;
mem[37] = 144'h0018fe9000a50108ff15fe08fe720086feca;
mem[38] = 144'hffa6ffecff7ffe7d0122ff4f0002febc00ca;
mem[39] = 144'hfdcdfe9dfe590131016501e1fe7f002dfebb;
mem[40] = 144'hfeef0060ffd3ff07016600f70004fdfefeb3;
mem[41] = 144'h0117feefff0e017d01df00acfe95004d0020;
mem[42] = 144'hff6dff7ffe08fedf014800c5012f018dff5e;
mem[43] = 144'h0082fef5ff0100420158009800f400e80160;
mem[44] = 144'h001501280037feddfe5afe3c01a000050100;
mem[45] = 144'hffd1fe41014a0037ff9cff350030fe4efff2;
mem[46] = 144'hfe8aff9ffe30fe14ff9dff82ff45ff800010;
mem[47] = 144'hfe48fdebff81ffaffe9cfe6300f2000e00ac;
mem[48] = 144'h00f6fff2fe22fdeeff94ffcdfda8ff4cff2c;
mem[49] = 144'hfe6700db0050fdb6ff1afe85ff5fff0f00f9;
mem[50] = 144'hfe27fed701c0011c0046fedbfda600b5006d;
mem[51] = 144'hfd830086fd8ffe32002bfddffed6fd79fee4;
mem[52] = 144'h000dfd6afd5dfd8bfe43003ffdde0050002d;
mem[53] = 144'h00cc00ff0092ffa100fcff06ff7c01340088;
mem[54] = 144'hfefbfea3fdaaffc8ffeefefdfe8eff26005c;
mem[55] = 144'h00b40030ffb1fe520062fe4b0101000ffee1;
mem[56] = 144'h0108feaefe59005a0029fed9fd83fefdfe10;
mem[57] = 144'hfd770097ff35010bfdd8fe34fd8f00a5ff90;
mem[58] = 144'h0007ff9d00e7fe4fffdfff6900f4ff7f008d;
mem[59] = 144'hfe71fd78ffb9ff5aff07fe77fd7cfeca00b9;
mem[60] = 144'hfede017ffe400054feb80144002b00f00120;
mem[61] = 144'h018400550071001a00ef00b90122fec7fedb;
mem[62] = 144'h0010fef3ff3afe2a0013ffa3000bfec40036;
mem[63] = 144'hfe2cfd54feda0083fe9afe29fe910108ff63;
mem[64] = 144'hfdc0fcaefe72fdc5feffffbffe4e00330247;
mem[65] = 144'hfdc6fa36ff6afce8fe20fd90ff4bffad0216;
mem[66] = 144'hfeb3fde60126fc2dff02ffa102fa04a4ff80;
mem[67] = 144'hfaf2fa5b01a7fd79fd7a022dff1c048b0260;
mem[68] = 144'hfcf7fc32024cfe7bfd4501a800c60132016a;
mem[69] = 144'h062dfd79fe6d0024057608c704b5015f0087;
mem[70] = 144'hf85200cb0201fe2ffe13ff3a00da0519fe5c;
mem[71] = 144'hfd280400041d01c0013cfd1cfc0f0302fede;
mem[72] = 144'hfeb8fcdf013aff38fdb6ff74ff4f0279043f;
mem[73] = 144'hfe4cfce2fef6fb52ffae0043006d032e047d;
mem[74] = 144'hfc9ffba3015bfea5feb7fd72fff2033904d3;
mem[75] = 144'hfef1069f02c5009f010a05c9092f06ebfe74;
mem[76] = 144'h0183fe3a00d3ff19fff70081ff5dff74ff4e;
mem[77] = 144'h0108ff4a0104ffe600bbff4cfe81000ffe47;
mem[78] = 144'h006dfbc9fe93fd87fefafcd5ffacffc40536;
mem[79] = 144'hff81fadbfe46fec1fe4e0136008902720367;
mem[80] = 144'h00fcff8efeffff77ffceffa4ffe7001f017c;
mem[81] = 144'h0178feb300f200a200defe8efea3ff9ffe54;
mem[82] = 144'hffc1ff30ff23fe0700a300a70120fee2007e;
mem[83] = 144'hff1d0008006e01180127014c00bb00a0fed4;
mem[84] = 144'hfe790158fde1fff7ff990127fde8fef0006d;
mem[85] = 144'h00f5008afdf7ff8000c80000ff12ff2b0034;
mem[86] = 144'hffc20000fdfafeb3016000f001caff0dfe92;
mem[87] = 144'h016301230234005201c8fe35fff901fcfe33;
mem[88] = 144'hfeb300c3fe240009fe51ff71013fff8f0020;
mem[89] = 144'h00c3ff620087ff98febbff98ffbafe5901b0;
mem[90] = 144'h00a0feb7001efe5300170050ff2d009a00fe;
mem[91] = 144'h011eff4cff69fe89feccfdc8ff390033fffd;
mem[92] = 144'h0151fe6ffef3ffc3019cff8001e1018a00c3;
mem[93] = 144'h00de014a00dcfec1ffb50196000f009effa9;
mem[94] = 144'hff3501740066009d001b007cff7efe2afe92;
mem[95] = 144'h0117feae00690092fe5a00220129ff7bfdc0;
mem[96] = 144'h041403c1032ffb29007901d002c40283049c;
mem[97] = 144'h0146014405f8fbcc0050047e038502e5058e;
mem[98] = 144'h00b804ad051cf9a1fa4df8d2f930fde7ff5e;
mem[99] = 144'h03da048807c80109ff42002f02d90241ff39;
mem[100] = 144'h034904c204a0fd2dfc790140015b012cff73;
mem[101] = 144'hfa740014ff66017ff8c2f3faf95dfef700ca;
mem[102] = 144'h041007a00558f9e1fa3dff7a01edfff400f5;
mem[103] = 144'h049d058e01d1fdbff99bf65bfc69fc36fe2f;
mem[104] = 144'h01ce021204a200b90071014a045d02270375;
mem[105] = 144'hfed90504063bfbcfff3000bb0157021b02a9;
mem[106] = 144'h02d504f007b2fc93fcb5ffad0142017501c4;
mem[107] = 144'hfb7efc3dfc31fecd0112fabbf4f6fa90fe47;
mem[108] = 144'h01e4fea40071feaf01c5000dfe6602400156;
mem[109] = 144'hff2e01acff70ff42000600af0142ff1bff89;
mem[110] = 144'hfefa017403c7034e01fc05e00256065c06c4;
mem[111] = 144'h011301860423000aff73002900d701b20586;
mem[112] = 144'h0086fec7fe65fe770138ff06ffa9fdedfeae;
mem[113] = 144'hff12015ffee20076ff89febefe2b009dffd6;
mem[114] = 144'hff1c00a9fec6feac0011002e00bc0045ffc4;
mem[115] = 144'hff2b012afdf80008fe9000c6fee1ff54fee8;
mem[116] = 144'hfe0e017300e4fed50100fe1effb4001aff65;
mem[117] = 144'h002c00a90171feadff65fe87000f013cff42;
mem[118] = 144'h0025fea4fe40fee2ff4efe06ff6900fafe45;
mem[119] = 144'hfee2fe67fe5ffdc3017a00e5fe8a0091feee;
mem[120] = 144'hfe400139feb9ff760016ff5dfe89fde2ff04;
mem[121] = 144'h00d8002900230176fe3d00e800b4fddcff0a;
mem[122] = 144'h007400a3007301e900ce0155fe89ffa8ff97;
mem[123] = 144'h009f0031fe58014cfeabfed8ff960213ff09;
mem[124] = 144'hfe4601c10153ff26006501b9fede01740159;
mem[125] = 144'hff8f001fffbcfe89fe51004a0048fe4a0122;
mem[126] = 144'hfff7ffb9004cffe4fdf101300055fe3000ca;
mem[127] = 144'h0128ff6dff2a0037016bfeb7ffd6ff250017;
mem[128] = 144'hfd46ff8cfbd8fec9ff61fed5005a0042fce1;
mem[129] = 144'hfd46007dfd8dff70ff2a018c0323fe0dfd7d;
mem[130] = 144'hffc9fca1fb0e02f2ff010255039c01d70179;
mem[131] = 144'hff6fff13fb7cffdbff3b03e10162ff74fcf6;
mem[132] = 144'h0075fff1fb95002b0261035201a3fea0fecb;
mem[133] = 144'h048801a900f600ad01fe0451054601a700c8;
mem[134] = 144'hfd50f98efccc0318fee4ff47feabfc720198;
mem[135] = 144'hff62f948fdb30416fea200aeffaf01d50249;
mem[136] = 144'h00a6fdaefdcbfd87ff9f029000effeb9fce2;
mem[137] = 144'h003ffd55fba9ffcb00ef01b402f1feb1fc8d;
mem[138] = 144'hfe07fd0afde2feb80307039e039e0111fe40;
mem[139] = 144'h02f4071c03be018301ac06bb02160267025c;
mem[140] = 144'h01d7fedbfeaafeafff8ffcea0019fff70199;
mem[141] = 144'hff7301d20192ff40fff3006e01540108ffa0;
mem[142] = 144'h0059feb2ff82fe65fbf8fe3b0175fff4fb11;
mem[143] = 144'h0000012cfc75fdc7fe280039038bff5efbde;
mem[144] = 144'hfcd801650438040c019f03fa00edfdc2fee7;
mem[145] = 144'hfdaa00ee02520479027800e600f8fdf001a8;
mem[146] = 144'h0423030eff8f018f02910899045f0043ff78;
mem[147] = 144'hffff0181017001bf02b500d90365014a0000;
mem[148] = 144'hfec4007c02d7026a0347011a02fa00b4fe19;
mem[149] = 144'hfde100f502a2ffe7002302c50349fe7f00d7;
mem[150] = 144'h01a5007c0196ff130254060d049c02090205;
mem[151] = 144'h07e2fee5fd48fff801fc071c077d02950111;
mem[152] = 144'h0162012e02b40463009c03c40213ffd6010e;
mem[153] = 144'hff0dffd0016e027403ef0145fe36fca4003e;
mem[154] = 144'hfe5f019d0438006a02d8038f01be0215001d;
mem[155] = 144'h05cb0083012c012bfcfcff74fe47032cffda;
mem[156] = 144'hfec6ff85017a01ddff24ff57fe29fe6900cf;
mem[157] = 144'h00a0ffc9ffd3ff2a014dffc9fe4bff52feb0;
mem[158] = 144'h0081038701da05280123014c00b7febd025f;
mem[159] = 144'hfe8b001d031c05cf029000bc0261ffbdff38;
mem[160] = 144'hffa3feb4ffc4ff990070ff24fadffd1f0079;
mem[161] = 144'h00f3ffde00d1fd4efe95ff2afd70fd6b00fa;
mem[162] = 144'h0177feb902fbffc006d0034500f1040b0414;
mem[163] = 144'h0232fa530179fdd2ff9402c2fdc2ff8c01f0;
mem[164] = 144'h0083fc39ff8e01c7ffd90240fe20fea90118;
mem[165] = 144'h0453010ffe8b0186ff96084c01f6fe16026f;
mem[166] = 144'hfd90fc49fecf012206ac044ffe4105da01da;
mem[167] = 144'hfcccfed001e6023807740934052e073402d4;
mem[168] = 144'h01e7ff0c00affe5a0092feecfe0efc6f0336;
mem[169] = 144'hfdec002b01f3027300b9ff00fbe2fc7d03b7;
mem[170] = 144'hfc60fbea00d6fe9c00fefe53fcfbfe0900d9;
mem[171] = 144'h03f102a5015fff2200fe03b3082b0d9903be;
mem[172] = 144'h0173ffd500d7ffbdfff8027aff2bfff800e0;
mem[173] = 144'hff990060ff97ff77fec8ffeb009c01a3ff5e;
mem[174] = 144'h032b01b00065ff31fe6dff95fda8fd2effa8;
mem[175] = 144'hffb8ff8bfee5fed6ffa5ff10fbdafcc80122;
mem[176] = 144'h012f00f9ff64fe7200fe00a2fffefde4ffd3;
mem[177] = 144'hfe18fe25febaff9a00d8febdfe31001300f2;
mem[178] = 144'h006901c4fee801d50015013afedaffd7ff26;
mem[179] = 144'hfe48fdc1009c00edfe20fe1cffe1fe9d0176;
mem[180] = 144'h00e501370066fe47fffd0139008fff36001a;
mem[181] = 144'h0169fedcfe8e011e00d500cf00a300ecff17;
mem[182] = 144'h009f0136006cfde5fee2fe99ffa6014fff6b;
mem[183] = 144'h017301000144fdfcfedafebe008f0052fecc;
mem[184] = 144'hff54ffacfdc8ffa4ff04010dfe85fe98fe6e;
mem[185] = 144'hfe180133fe11fe24023f0070fe8401daff2d;
mem[186] = 144'hfee7005500a90012007800f4ff00ff120030;
mem[187] = 144'h0158014500fa0048fec4fefaff28fec9ff2d;
mem[188] = 144'hff52008a011fffbaff320080fff8fe4600a9;
mem[189] = 144'h01690074ffda01a4ff18012d01bffe32017c;
mem[190] = 144'hff11ff9efe47fe23feedfe63fe74ffb500c9;
mem[191] = 144'hff0dfef6ff4e00ccfe54ffadfea60166ffc5;
mem[192] = 144'h027000e6ffc0fdf5016eff810277fea1fdcb;
mem[193] = 144'h0300024e00cafe2500940205019cffaafd60;
mem[194] = 144'hfd7efbaffe330198fdfafcb0fc1dfd31009d;
mem[195] = 144'h00abfdcefe37fe27fedf0111ff83ff0efde0;
mem[196] = 144'hfebb012ffff5fe53011e004702adfd72ff95;
mem[197] = 144'h0021fe14ff3dff9800f4fbd0001a002bfd47;
mem[198] = 144'hfe950044019bfd1afbe3fe82fc7afdf2005a;
mem[199] = 144'hf819fd0cffa2ff52fbd6f998f5f3fca3fe4f;
mem[200] = 144'h00af0194ff78fde8fe1f0210029800b2ff94;
mem[201] = 144'hffd3025a017dfd65006202800349ffc4fe6e;
mem[202] = 144'h00a7020100a0ff0d010000bfff4f0043ff7a;
mem[203] = 144'hfbd6fc43feb4012f014b0210ff71fbdcfe38;
mem[204] = 144'h0263ff40011700e700d5fdd3ff270207febd;
mem[205] = 144'hfefaff1c00bd012eff1e0052fe6afe8f010d;
mem[206] = 144'h02d201510120fdf300a30258019b01d2fe2e;
mem[207] = 144'h00cd00cb0077fdfbfe0f0177005efea10021;
mem[208] = 144'hfe1dfaa6face03280224fddffe18ff81fd3e;
mem[209] = 144'hfdb3fb1afc5c04ba00e4fbf9fd50ff190045;
mem[210] = 144'hff03f9cc0171092b065d0461084801f40219;
mem[211] = 144'hfdedfc14fcb301ab01e9013bfbe301a001c2;
mem[212] = 144'hff85fafcffbd027204520197ffe402c50283;
mem[213] = 144'h079700d4ff60011f0b110f8904480493007b;
mem[214] = 144'hf9affd10002404ea09b2ff52fc3b0339027c;
mem[215] = 144'hfa8403050224031b08e708e8045b027e0122;
mem[216] = 144'hfd8efcfefbef0236032cfe78fd29ffc80086;
mem[217] = 144'h01a5f9fbfe25049802c1fe3aff6201710274;
mem[218] = 144'hfcc0fc10fae105b70389fdd7fcf803e40360;
mem[219] = 144'h07fd06e901fe0237013508f7154609ae001b;
mem[220] = 144'h017d004c01150016ff44ff6c02c4fe6d002c;
mem[221] = 144'h00200000fe96ff01014000f900f6fec9ffba;
mem[222] = 144'h016efd15fb81fdc7fc76fc2ffd94fd7ffe59;
mem[223] = 144'h004bfd1efd4c0219ffeefe9ffdf1016701d6;
mem[224] = 144'hff76feff0012ff3e00f0023a0258fee403ed;
mem[225] = 144'h000801e0ffd5feeb01170333031dff4e0153;
mem[226] = 144'h02de016f026cfe2903d905b6022701eefeeb;
mem[227] = 144'hfe9efd890337004ffdd601e003d10415021e;
mem[228] = 144'hfe9601540108fe3800280272018e020a01ba;
mem[229] = 144'hfcf5007bfdf5fee4fcfafc8803cd00d6fff8;
mem[230] = 144'hfe2001ce0357fc8a023a06e002e601dfff3f;
mem[231] = 144'h05cd00e2026bff69004c0297037702ddff0f;
mem[232] = 144'hfd53ff5301aa015f00e0016c00000265015c;
mem[233] = 144'hfe090069025afec7013e0320fff8fd4d0198;
mem[234] = 144'h0115ff7104dfffb2025a06020320035a027a;
mem[235] = 144'h0273ff3b000d00f9003afddbff4601af00bb;
mem[236] = 144'h007401dd015101610138011bfd89ffd20068;
mem[237] = 144'hfecafee70189006d00c60026ffe4002cfecb;
mem[238] = 144'hfe0d004cfdc1008600e6feb3fd78fe3f03f8;
mem[239] = 144'hfe10ff38034a008e005f01ad0161007b00ef;
mem[240] = 144'hff3f01d00197ff12ffe800d00180008d004f;
mem[241] = 144'h02fb003ffeaffe790039022501f00146ff37;
mem[242] = 144'h04130104fda8fe0efe5ffd31ff9d010b002f;
mem[243] = 144'h03220141fdda008f014701dc02f4ff590198;
mem[244] = 144'h03a1004a010fff52fedd01e9011d01d201f4;
mem[245] = 144'h028404bd00dd03a3fb3efd4b0210004b0364;
mem[246] = 144'h034ffb0cfb33025701adff32ff5affad00b4;
mem[247] = 144'h01eefe6a0062ffe202b4fc39fec9032803ee;
mem[248] = 144'h02ad002c0097fe1dfede013401ae02f5ff38;
mem[249] = 144'h0031fd4cfdf9008cff24019f0208ff6d009a;
mem[250] = 144'h03e20119ff38ffcf00c1ff2bffdf0100fe9d;
mem[251] = 144'h02df06d103c9ffa301780259fc51017503e0;
mem[252] = 144'hffb9005000f90017fed6021f018eff5afec9;
mem[253] = 144'hfe2ffe51ff30014300aefec4fedefe86ff8c;
mem[254] = 144'hff50028a0049fe410074043a0297028e0192;
mem[255] = 144'h013e020600b700bdff8e0285019301600257;
mem[256] = 144'h023803ec027d004e000003c4041402d500ae;
mem[257] = 144'h01b6052a02d3ffc20070043c044903affdbd;
mem[258] = 144'h02170277f86bfc08fbae00cdfd670124fded;
mem[259] = 144'h040203c00087fd9afdfb008e02aefe87fd59;
mem[260] = 144'h02cc062cfe86fe45005e03430197009bfe49;
mem[261] = 144'hfbc204f3015bfffaf7a8f2b4ff89fe5c00cb;
mem[262] = 144'h04c9fdf9fe52fd24ffa004160139fd86fe36;
mem[263] = 144'h0440f7e2fc1d0003fe19ffbfffc3fce7021e;
mem[264] = 144'h02f505f10149fdd90070044e02710076fe86;
mem[265] = 144'h0170069701e600a0018901c2003affa4ff15;
mem[266] = 144'h04a8034dfffa004a0052035402cafe55fb42;
mem[267] = 144'h0262ffe2fed5fe8f012cf998f4fffb2e021f;
mem[268] = 144'hfeb0fd78fd5d00ccfe910033fd41ffee0171;
mem[269] = 144'hff3400ef013a009c009bff4c00fd016b0128;
mem[270] = 144'h00ef02a701a40063024101cb04050316ffb3;
mem[271] = 144'h044404620360ffbefe7c02b602bb0179ffb8;
mem[272] = 144'h03b704c70415fb3bfd6e012f006301a704b7;
mem[273] = 144'h02d601a504c2fc40ffe4009a013000610369;
mem[274] = 144'h006f062406dbf85bfbccfcbdfaa301a4fe69;
mem[275] = 144'h05a204bc04e7fd73fdd8fdf3fec401200130;
mem[276] = 144'h00d303300209fd31fc91fd55ffad0002ff65;
mem[277] = 144'hff150081fff1ff38f811f3cdfac8fc900248;
mem[278] = 144'h05a2024a0347fd40fc3bffa7014e0020ffec;
mem[279] = 144'h047e02a70369fea9fc32fa5affe701cafdee;
mem[280] = 144'h037d01e502fbff15fe650205fe8900320266;
mem[281] = 144'hfe8e00510371fdbdfe01fdc1ffe0fd6d02b2;
mem[282] = 144'h016601ac028efc37f9cffce8fe63fd0dff4b;
mem[283] = 144'hfb17fe310163fff90157f7b4f485008cff4f;
mem[284] = 144'h006bfe50006bff700118ff6cfe7fff96ffbc;
mem[285] = 144'h0067001d00d3007aff46ffc5ff28ff3dfe1f;
mem[286] = 144'h00c5040900ad00d8026805810193014a031f;
mem[287] = 144'h01fc01ad01ddfdab00570095001900af0150;
mem[288] = 144'hfebf004301f9ff47014dffe500dc032700be;
mem[289] = 144'hfe8affaa006a017a01a7002d010102a7028f;
mem[290] = 144'h00fd0076fca8ffb90177076a062c06b8fe7c;
mem[291] = 144'hff8cfffc02b7fe7efff503e403de02d8001e;
mem[292] = 144'h00a10280008401dfffe002f103a802c4ff24;
mem[293] = 144'h004a044b02ad0019fd32fe1a01b6016301fd;
mem[294] = 144'hff84fc9bfdf1fecc03d506c402c7fdd600d4;
mem[295] = 144'hfe0afb15fd49ffe50290060303deff7d0094;
mem[296] = 144'h00db00af007efff4018100ca0267042800c0;
mem[297] = 144'hfeab014b003601b1025300f3023900f0007b;
mem[298] = 144'hfd3701ad02fd0042ffcd04dc020200dc0113;
mem[299] = 144'h04c00ccb04a7ff76ff65fe34034306c702de;
mem[300] = 144'h00f1ff150152fff20108fefe009d01a7ffb2;
mem[301] = 144'hfe7f00acfea5ff4efe65fe9fff76000001c4;
mem[302] = 144'hfdadffb2fdcf02c8ffacffdbff1400a50350;
mem[303] = 144'hfd9d02d1027d00c2ff1900f4006f00c602c4;
mem[304] = 144'hfd97feacff5afe5dffe7003eff180056fe72;
mem[305] = 144'hff81fdd700c7fe1eff7aff0bfdd9fdebfdd7;
mem[306] = 144'h013b010c004cfe1ffe16fea900bdff49fe14;
mem[307] = 144'hfde1013ffff2ff75012c007a0148ff45fe80;
mem[308] = 144'hff46fe280168015afe72fec6ff71ff2a00d9;
mem[309] = 144'hffd20045fe42fe84fda3ff2efed9fe5cffaf;
mem[310] = 144'h00a6ff77000efe9cfdb7ffcc0082fe64016e;
mem[311] = 144'h00bd005300db00e4fdf1ff76ff9fffeeffce;
mem[312] = 144'h01460108011d00f5ff0afee40067002e00de;
mem[313] = 144'hffd700e1fe21010b0117fe9cfdc40107fdd8;
mem[314] = 144'hfdb4007cff00fddbfe290155ff70fe620095;
mem[315] = 144'h0036005cfefcff8eff36005fff8200be0112;
mem[316] = 144'h011d0057ffabfeb100ad0191000800320071;
mem[317] = 144'hffe5fe6effbf0048fe630012fe4cfe8f0164;
mem[318] = 144'h013efef00129ffc2ffd2fed4ffc6ffeeff56;
mem[319] = 144'hfde2ffa8015fffa6ff4bfec1ff720071ff1a;
mem[320] = 144'hffbafef7fe390265005cfc23fde9ff2ffbbf;
mem[321] = 144'h01d30060fc8a02030009fdafff7c00a6fdd3;
mem[322] = 144'h01a2fbe5fdb6050a0315023500ceffea02a7;
mem[323] = 144'h0271feb1fa0302180335ff30fbf6fd4f02fc;
mem[324] = 144'h022e00f2fc3503fc020300850057fece020d;
mem[325] = 144'h022102f9fedf019706570a72027301e0ff7a;
mem[326] = 144'hfe64fa67fc3303a406c50065fca0ffe401b1;
mem[327] = 144'hfe95fd6300b104170658083efdef01ec0102;
mem[328] = 144'h0265fe52fbd0013f0201ff43ffdf00e800ac;
mem[329] = 144'hffaafec6fb4b05d0fe93fdb8ff80ff6fffb1;
mem[330] = 144'h00e0ffc9fb2802800330fe7dfdfafe5001ec;
mem[331] = 144'h05a600bd025b0092013a06b60ae403ac030b;
mem[332] = 144'h005eff90ff480159006ffd9dff57fcdc0059;
mem[333] = 144'hffdefe46ff40fe83016900ac0110febafeae;
mem[334] = 144'h00c2ffd0fc7bffe4fcd401100025ff87fbcf;
mem[335] = 144'h021aff98fc3f012fff0000d9ff230037fd39;
mem[336] = 144'hffbd0030fe09fbe7fcdd004c01d8ff5bfc48;
mem[337] = 144'h0181ff66fdb4fb6cfd0700c4031f0203fdab;
mem[338] = 144'h0074fbfbfba9ffb4fd4fffec0251ff52ffe1;
mem[339] = 144'hfed5fe58fba8feb4fdb600c403e3fea5fc5d;
mem[340] = 144'h01170164fd330121fef7feec033eff7bfd47;
mem[341] = 144'h0393021d017c03bc0145fde7037403bdff39;
mem[342] = 144'hfbf8fce2fc69009dfff4feaaff2aff8fffa5;
mem[343] = 144'hfdd8fb0dfe1301b8fd94fe1afc94000700a3;
mem[344] = 144'h0136fe54fef9fd02fe2600fe02f00006fe17;
mem[345] = 144'hfff90157fef1fee5fd30024b02b200c0fd11;
mem[346] = 144'hff26fea1fc72ff9cfdb8ff7b02f9ffe2fdec;
mem[347] = 144'h007903ad0047fcb3fe9704b701b1ffdc0227;
mem[348] = 144'h015dff43fe04ff550038fee6fee00108018e;
mem[349] = 144'h009cff7401030157023100a7ffb200fa0193;
mem[350] = 144'h0241fef4fd29fb8dfde6fefb00720027fe51;
mem[351] = 144'h0191ffb0fca7fe76fc33009403130038ff1c;
mem[352] = 144'h012e02010234fee3ff1dfbb6fe78fd5e0044;
mem[353] = 144'hff63015103e7ff87fe49fbbdfd86ffe20254;
mem[354] = 144'hfd35fd6203e0fc27fd9efa56ffadfb0dff83;
mem[355] = 144'hfde8010f023a000eff96fbd7fd2c00de00c8;
mem[356] = 144'hffd301bb00e90135fd3bfdcefd910166fe11;
mem[357] = 144'hfe5b0085fe4bfe8e03670814fd2001f0feaa;
mem[358] = 144'hffcd011901d3fea1fcf0f9e0ff820029ffd0;
mem[359] = 144'hfeaa030902d6fdbfff6100a0048301310039;
mem[360] = 144'hfff10172038f00c4feacfc5efed70064ff22;
mem[361] = 144'h0016016800cdffd7fed1fbc6fdf8028d0187;
mem[362] = 144'hfde2ffe9001eff68fdf8f9b3fd99ffdcffe5;
mem[363] = 144'h0180fc0ffc88012dfdbeffc707d9017a001a;
mem[364] = 144'hfe8a0167ffa3005c0226ffe1fe5e00610081;
mem[365] = 144'hfe55fefbff25ffd40152fe6f01d3ffcbffc2;
mem[366] = 144'h010e011502b101a002ebffd7fe6800f302bc;
mem[367] = 144'h00a500b00135ff4affebfcc3fb69010ffef5;
mem[368] = 144'hfe75fdcf006c00ec00ee00c901c1fe4e00a2;
mem[369] = 144'hffc4ff1effbbff2bfe65ffe8ffaffe00016c;
mem[370] = 144'hfe58ffc301db000eff5c01c501970041fe57;
mem[371] = 144'hfeb6ffda00cd00fa003800befe16ff4afdc4;
mem[372] = 144'hfe35ff3a004c0103ff26fe10fe99fecfff09;
mem[373] = 144'h005f0021015700d1fe2fffe1010800ccffe7;
mem[374] = 144'h00c5011fff4a0112ff86016300d8008bfe35;
mem[375] = 144'h011f01e1ffd9008affa9fe240178003e001e;
mem[376] = 144'h00040045fffbfdd6fee8ff2afeb5ff41014e;
mem[377] = 144'hff800166ffde0083014cff92ff47007aff86;
mem[378] = 144'h01b600d50003fff101c001c100d1ffcf0163;
mem[379] = 144'hff02003500870027ff62ff7000defea70107;
mem[380] = 144'hffc100880033ff4701d6fe4bfef001d4ffc3;
mem[381] = 144'hffad006bfe5eff32013eff98fe6301cdff1a;
mem[382] = 144'hffd70124fdcc009dfed10091feb000c200b2;
mem[383] = 144'h00ef009100dcfe7dff01014bff2b00bafe29;
mem[384] = 144'hff4eff10fe10ffdafecdffa7ff74ff65fe0e;
mem[385] = 144'hffd10052ff8a002bff57006aff6000af019c;
mem[386] = 144'hffdbfdbffeba00160115fef2002cff9c008f;
mem[387] = 144'hfddf0177feabfe6bfd7f0056febe0090024c;
mem[388] = 144'h0029ff19fd94007affaefd2ffe32fff101a5;
mem[389] = 144'hfeb8fdb30044014bfecdfe930070fff2fff6;
mem[390] = 144'hff49ff6dfd94fdac01de0023ff66fe6400ed;
mem[391] = 144'h00f5fffaff85010d011300e8ff55ff630074;
mem[392] = 144'hfdebfeedfee4008c0036fd8a00eb0060fe48;
mem[393] = 144'hfe8700a4fdc8ffd9fd98fe5cfdd9ffb8ff99;
mem[394] = 144'hff2b008b0003fec0ff31fd52002e0019ffae;
mem[395] = 144'h029cff29fe60fe1fff8cfd7b0290ffe500ef;
mem[396] = 144'hff1001d7003a016d00d9002dffbfffe3fe4c;
mem[397] = 144'h010b0037ff83feda01cafef1ff4700d40088;
mem[398] = 144'hfeeefeb0fe1efea90073ff61feebfe01fefa;
mem[399] = 144'hffbb0166fe31ff77005900570059fe580130;
mem[400] = 144'h0044feb70023ff25feb2f92ef998fd44000b;
mem[401] = 144'h011eff1dff57feeefe60faf2f935fc61010d;
mem[402] = 144'hffa0fa9e035601c502b203be068600970355;
mem[403] = 144'hfc04f9eb02c7fecffe34fac2fbffff42022e;
mem[404] = 144'hfcedfade01f00362ff0dfdc3fe2401350262;
mem[405] = 144'h03ebfd64fe2102c809480ca200fc00ef00c2;
mem[406] = 144'hfacffd8c030d03da052bfdd2fd21040e031d;
mem[407] = 144'hf752021f045e042106b50c58070d0548ff5f;
mem[408] = 144'hfdb7fcef00e2ff80fcdafacbfa99febf01bc;
mem[409] = 144'hff8bff380158032efc80f8c5feb0feed0121;
mem[410] = 144'hfba8fd1bfecc0165014bfb11fb5201200324;
mem[411] = 144'h0790015402adfe66fdbf036a1060096e021c;
mem[412] = 144'h01380222ffdb017dfefdfff1ff2b0038feb6;
mem[413] = 144'h0118fe96fff70022ff7100d60012ff08fe2c;
mem[414] = 144'h01dafe6102440059fedbfb4cfa34fe39011e;
mem[415] = 144'hfdfffdf9fec8ff41ff36fcacfadcfd530040;
mem[416] = 144'hfbc2feb7fc91fd52fce40025ff78ffc9fe2c;
mem[417] = 144'hfb4bfe65fe22feb2ffafffcc00c4ff4cff74;
mem[418] = 144'h00d30150ff97fe1202610171ff50fff501b8;
mem[419] = 144'hfd96fdcbfd27ff15017c0265011f013efcb8;
mem[420] = 144'hfdf2fda6fea70273fde00117007bfffeff65;
mem[421] = 144'hfd33ffc80051fdabfd36ffaffd74ffa4fe22;
mem[422] = 144'hffc2ff22fb8101fc017b02e001b1fec0fd46;
mem[423] = 144'hff62ff17fd1cffd5ff84ffa3ffaeff4efe6a;
mem[424] = 144'hfbe3fe61ffccff60fd3301e8ff0c00df0015;
mem[425] = 144'hfbf6fe43fcfcff70fe6001f3019dff630013;
mem[426] = 144'hfe3afd69fd39ffe5fef0023c008a0178fc32;
mem[427] = 144'h00a1008efe45fc5900d6003bfeafff1afe98;
mem[428] = 144'h00c8fe58feb501c5ffd9fe9fff0bfefc0156;
mem[429] = 144'h0069ff82fe2f011b003afefdfecf010cfe47;
mem[430] = 144'hfd88feb2fe19fb22fe97fdd6fd38ff11fd41;
mem[431] = 144'hfdb8fd72fcccff58ffa8ff62ff720028fdd5;
mem[432] = 144'hfe88ffc0fe160066012effa10035fe1f0017;
mem[433] = 144'hff41feb40113ff8c012aff71fdd7fe92fe1b;
mem[434] = 144'hfeb10174ff66feab015ffe50fe91004d000d;
mem[435] = 144'hfe4c0122fe020101ff02fe6efed9007cff5c;
mem[436] = 144'h0062fe2d003c0084ff59ff81000400c800ff;
mem[437] = 144'h0034ff1bffe80155ffbffdce0009fece0160;
mem[438] = 144'hfea3ffd60129006100c9ff17fdf0ff2f0046;
mem[439] = 144'hff41fe7b007800c4ff020089fe1100cc0113;
mem[440] = 144'h0137ffa600aeff8dfe1c013dff9b0027fde0;
mem[441] = 144'hfdd4018e00390023002afed5ffd501cbff5b;
mem[442] = 144'h017a0015ffed004f0035ff30fe83fef6012a;
mem[443] = 144'h012cff1e011fff57fee2013bff9500c0ff22;
mem[444] = 144'h012e0107ffff0061003fff56004c00f7fea8;
mem[445] = 144'hff9900370093ffdf0171ff9300ff00baff50;
mem[446] = 144'hfe65fe04ff8afdc1fe49001300c9ff3300eb;
mem[447] = 144'hffc50158fe6a013b01740134feebffc20000;
mem[448] = 144'h0061009400460043feaeffedfde9fe640175;
mem[449] = 144'hfe3bffac009700d40149ffe4ff96ff55009c;
mem[450] = 144'hfe4dfe5001a2002eff14ff64fe47fe6fff8c;
mem[451] = 144'hfdc3fe94016500d700cd010cfe910068ff4c;
mem[452] = 144'h0121ff04ff42feb4fe22fec1ffb0000cfe9c;
mem[453] = 144'hff840012fec9001900d6ff4700710010fe46;
mem[454] = 144'hff8ffdbc000cfee2fef300c5fffa01080025;
mem[455] = 144'hfeb3fe41003a0030ff4200f7fe9fffda00b1;
mem[456] = 144'hfe1500f8fdcf0088fe3bff37ff2900fffffd;
mem[457] = 144'h0070003a009affbdfe12010afe90fe590089;
mem[458] = 144'hfebbff55ffd900be006dff21ff7cfe61018e;
mem[459] = 144'h00840105ffc2ff28fec50074ff33010101fc;
mem[460] = 144'hff9b00f6010900420163fe5f0093feda00a6;
mem[461] = 144'h01aefe81fe4101c5ffe5016ffe75ff7800e4;
mem[462] = 144'h00690087ffbcfecdff8effde00dd00d100bc;
mem[463] = 144'h00e8015f00f0ff4efeedff24ff740035fdde;
mem[464] = 144'h034b01a7ff98fd03fe710005ff52fc9efdac;
mem[465] = 144'h0152ffd2ff89ff4e00b6fff700dbffa3fdfc;
mem[466] = 144'hfc3dfc8d0149009cff560022f92efa6e0054;
mem[467] = 144'hfe3aff3b0262fdc50097fe07ff2ffc1e001a;
mem[468] = 144'h016bfff3fef1fe95018f008efdf3fcaafd71;
mem[469] = 144'h0018ff63fdfbfef2ff3cfe88006cfd81fd0c;
mem[470] = 144'hfe0b0350017efe8efe22fcb700bf018efe30;
mem[471] = 144'hfb10006600e500deff6af683faa7fe4aff68;
mem[472] = 144'h02a60023007a004cfeedfeaa00a4fd3600de;
mem[473] = 144'hff78ff0cffcffecafd8d0128fe3ffd480065;
mem[474] = 144'h003e00bcffaffd02ff56ff5d0140fff7fe7a;
mem[475] = 144'hf5edf652fb800242002900e2f68bfbdefca8;
mem[476] = 144'hffdcff24ff9b0029fe42fe32fedcff55fe8a;
mem[477] = 144'hff74014301bdfef5ff4c0036ff88015bfefc;
mem[478] = 144'h0174003a0200ffb30095ff61fedafe2afeee;
mem[479] = 144'h018dfe490231ff5fffb8ff85feb0fcf20069;
mem[480] = 144'h031dfcc3fe0cffcd003e018602db030d0235;
mem[481] = 144'h0294ff7a00dbfeca0079fe41ffdb02ef0250;
mem[482] = 144'hfaa3fe2102800064fe89fc62fca6fb84ff71;
mem[483] = 144'hfcad02430302033b0384003801f304350329;
mem[484] = 144'hfda0020f017602dfff4aff6d03950185004b;
mem[485] = 144'h020a00f70081036307570329fdb402d901e0;
mem[486] = 144'hfdf208cb02c70204fb99fc1a05b1fd920038;
mem[487] = 144'hfc07057401ab01effe56f907fd03fab3fe1f;
mem[488] = 144'hff2fff9c01de021a0043006100c3005f0257;
mem[489] = 144'h008cfd730280febefd5a00fe026c040a01bf;
mem[490] = 144'h00540037001f019cff3cfd08000501fa0287;
mem[491] = 144'hfbefff7aff4500dc0237056001b8f9f50046;
mem[492] = 144'h00b400a500fcff12ffc8ffc600220123012e;
mem[493] = 144'h0131014a01a30158fdfc003000edfedb0149;
mem[494] = 144'hfdf0fb5402d1009fff9aff72029d048f013a;
mem[495] = 144'h007afcb70233ff8901b101420166fffe033d;
mem[496] = 144'hfd980104fe1bff2dffd1fe67fde6fecfffed;
mem[497] = 144'hff5d0017fed4ff200074ff66fe3dfdfb0104;
mem[498] = 144'hff0f009b00a2fe6c009e00a3ffd2fe3c01bb;
mem[499] = 144'hfdb200d700c100e5fe73ff7c00dfffe4fe0a;
mem[500] = 144'h00e2014e00f3ff29fffeff1afdb6fe2efdad;
mem[501] = 144'hff520109fddafe45ffdb0087fe2c009f004b;
mem[502] = 144'h001afe16fea100bffeebfff4ff9afe71fe72;
mem[503] = 144'hfef7fe7100d70120feb5011bff04ff7dfdd9;
mem[504] = 144'h00c200120020010eff3c00d1ffd9fe1b0024;
mem[505] = 144'hfdb2fe58fdce010301d401c4fe6400d5fdd4;
mem[506] = 144'hfef1fea700f8ff760094009cff1cffa900be;
mem[507] = 144'h0204ffd30104ffda00b7006d014e0101feca;
mem[508] = 144'h0061002efe3b00cf00c4ff25ff48fe280021;
mem[509] = 144'hfe8bfe7cff230099ffce00f6012cff8300b5;
mem[510] = 144'h00ecff7900cf006f0159fea0ff510149fdbd;
mem[511] = 144'hfe0ffec10158fea0ff310056ff10ffb4ffb1;
mem[512] = 144'h0030fe92ff49fa16faa7fcd6017e017b0073;
mem[513] = 144'h010cffbafd8afdd6fc22feed019d006f0123;
mem[514] = 144'hfd6efe2d00fbfd05ff68ffa60276fea7ff5b;
mem[515] = 144'hfdbefdb902dbfd5cff37fd4f0053041803db;
mem[516] = 144'h00cd010d012cffbbfd56fd89025f03ea00f0;
mem[517] = 144'h00d7010effba035404090369003105c7fff0;
mem[518] = 144'hfef606210448007ef9f7fded055b03d1ff95;
mem[519] = 144'hfc50036b041e0274002dfeb402f9fd9cff8b;
mem[520] = 144'hfe4bfe3b0069fbe4febafcec02970391ff62;
mem[521] = 144'hffa1ff0dfe79fda9fbf2ff700173040900c5;
mem[522] = 144'hfd6701a60038fd5dfaa0fd65020c05ec040a;
mem[523] = 144'hfd10fd5bfe69feae015b04ce0699fecdfedf;
mem[524] = 144'hfd9affc8013cfe28fc98ff63026f02ac013d;
mem[525] = 144'hffb7ffe2019cfe4d003600a200f601cfff6b;
mem[526] = 144'h005b0026ff4bfae5fe8dff0afeb900f1ffd8;
mem[527] = 144'hfee800dcfefffbc1feeefd77ff5701bfff88;
mem[528] = 144'hfca6ffae0185fee1011902960138ffff0181;
mem[529] = 144'hfcbefd92003f013c005102a6ffaa0068025b;
mem[530] = 144'h009c00b1ffea011301b2079909880959fe30;
mem[531] = 144'hfbc6feda03a9feebff2a02d5050c034d02ef;
mem[532] = 144'hfd01fe1c0211016a01d6040103d304310310;
mem[533] = 144'h015a01da02cf00ec01970241047c01230167;
mem[534] = 144'hfcdf01260108ff3502b5079f07e4057b02a5;
mem[535] = 144'h0051feab011b00c501870743078705e60273;
mem[536] = 144'hffddfdd2ff40ff830123001e030f032801fb;
mem[537] = 144'hfe14ff5cff8f003601ce032f0113ff5b013e;
mem[538] = 144'hfd0701490000fe5e000001d202cb0312029f;
mem[539] = 144'h0407092d07e3fffe00ad037d042b09c30099;
mem[540] = 144'hfeefff03fec6fe190058027f008a0226fec2;
mem[541] = 144'h0064fffdfe57ffab0051ffb8ff98010dfff3;
mem[542] = 144'hfee1fe20feba004e016afcdbfefd0175027f;
mem[543] = 144'hfc8efe6a0000fdc7ffa2027802e9008902d6;
mem[544] = 144'hffeb003c0013fdb1fdebfe06feea00780139;
mem[545] = 144'hff430137009a011efe44ff910104007c00da;
mem[546] = 144'h0013ff1a017e00f500dbfe9400c8ff6efea6;
mem[547] = 144'hff1d013efe79ffa9ff4bff0cffc1ff3fff6d;
mem[548] = 144'hfedc0011fdf0fdbafe56ff68ff61fe360120;
mem[549] = 144'hfdc6fef2009dfe000144feeffe3ffdb60143;
mem[550] = 144'hfe55ff7d00590027015bff97fe37ff38ff5a;
mem[551] = 144'hfde0003401b7ff5bff9d0114fe800120ff50;
mem[552] = 144'hff35ff33ff1effb4feb2fe0c0108009f00a8;
mem[553] = 144'hfe0b007ffdffffc1007afe75ff90ffbdff1c;
mem[554] = 144'hfe33feed0023ff7cff7cff56fe46fe3afe44;
mem[555] = 144'hffe4ff480077ff4c0006fddafe58016ffe35;
mem[556] = 144'h00d5012cfff800cbfe93ff24fe6d010bfe93;
mem[557] = 144'hfe44ff21ffaaff480168febbff5801750053;
mem[558] = 144'hff36007c0100fec9013effedfe85ff8a002e;
mem[559] = 144'hfea3ffb5ffeafe9d001600bdff73ff0cfe32;
mem[560] = 144'hfe44ffba00d4041004d3032c0123ff0c000e;
mem[561] = 144'hfe62021700ec0205035f04620166ff7fff3c;
mem[562] = 144'h05f20227f94c04ce069d077704be05570053;
mem[563] = 144'h02bf0211feb1027a02df027d01e1ff56ff36;
mem[564] = 144'h00f101c4ff16007101b2056803c60043ff0b;
mem[565] = 144'hf8300305021cfc62fca8fdcb03f0ff6f01e0;
mem[566] = 144'h02c4fb37fc9a017206a808dc03d8fef3019f;
mem[567] = 144'h05fcf845fd67006b0390062706cfff6bff74;
mem[568] = 144'hfe1d0101ff3f02fb0294047e0190fefa00a8;
mem[569] = 144'hfe1f003ffff303be0402023e008dfc34ff16;
mem[570] = 144'hfe71025a00f002a402c304680186fedefef5;
mem[571] = 144'h051c0774027e02b1ffc6fc4bfd8a046f0179;
mem[572] = 144'hfe3bff40ff57ff32010f0002ff34fdd80054;
mem[573] = 144'hfe8500ebfed8fe98017dfe9600dafe3c017a;
mem[574] = 144'hfe6e03cc00d203a601e5014101cafe26ff61;
mem[575] = 144'hff3b02effed302fd01d9047e01050200ffc6;
mem[576] = 144'hfe8101d202280253042d03960397ff74ffe7;
mem[577] = 144'hfd2e014c00eaffae03bb03e30417fef9fe9b;
mem[578] = 144'hfff3febefc5702990191064b018efe58fd0a;
mem[579] = 144'h0165008cfeb90049ff5704a70396fd4aff20;
mem[580] = 144'h0168fdd6ff62fe77028902de022dfd12fe4e;
mem[581] = 144'hfad3002efe11fd32fc85fdf605f6fdc9fda9;
mem[582] = 144'h0001fd41fe73fd96ff3803adfec5ff2afe79;
mem[583] = 144'h0237f693fc560057fdfc00befd85feb00014;
mem[584] = 144'hff02016aff420199011502d4005a002afe23;
mem[585] = 144'hfefb0162ff46fce601980296feaffe73ff20;
mem[586] = 144'hfdce001200abfdb301f60675048affc6ff30;
mem[587] = 144'h0053fdbaff5a025dfebbffcdfc62feacffcc;
mem[588] = 144'h0093ff0bfed40004fef40062016dffca00ed;
mem[589] = 144'hfe43fe8d000fffd3ff9cfe86ff0501400028;
mem[590] = 144'hfc810253ff7cff12007e0269029efd1fff4d;
mem[591] = 144'hfeca010effe4022f017a01e4034a00dbfe02;
mem[592] = 144'h002bfee1008d01faffaefe64010d00e1ff70;
mem[593] = 144'hff1efeb9fdc60073febdff42015ffec2fe8a;
mem[594] = 144'h002800e900b50041fdce01300050016efed1;
mem[595] = 144'h014e0110ffbbffc20028003700dc00e4ff8d;
mem[596] = 144'hfdfa003dfe990027fe08fdc7fdf300fc00a9;
mem[597] = 144'hffbdfdecfe6600e000d5013e0063fdf7feb1;
mem[598] = 144'hfdcfff8bfe1f00c1013cff16fef0ffb2ff26;
mem[599] = 144'hfe51fe8701520065fe3600460044000fff94;
mem[600] = 144'h0090008f009700ebfedbffbdfee3fe68fdf4;
mem[601] = 144'hff50fea8ff52fdc3ff4a0147fed7ffcbfeab;
mem[602] = 144'hff28fed100bafeec009e004200deff92ff46;
mem[603] = 144'hfe26ff370031fff3fe610042ffa0fe6b00d9;
mem[604] = 144'h01970056012401c500980194ff16000e01b7;
mem[605] = 144'h0183ffcf0074017000cbff2bfee201a900e0;
mem[606] = 144'h0072ffc700c5fefcffc0fe33fea4ff560129;
mem[607] = 144'h009400f20095ff59fe73fe8b012f0029001b;
mem[608] = 144'h00a30097021502b8fe4a000401ed00470370;
mem[609] = 144'h001efed301dd030400a50022ff0200b00295;
mem[610] = 144'h005801320530fff900e20521053d040b01e9;
mem[611] = 144'hfed00000015f01fb0028020d03a103cc01fd;
mem[612] = 144'hfebf004400a701d9027002710334017b022d;
mem[613] = 144'hfe9a039800370183fceffe25fe4501ae00ef;
mem[614] = 144'h005e005f0122011d06a706cb045d06b40208;
mem[615] = 144'h0224048c03a2007f06710b13096605a503d1;
mem[616] = 144'h008d01a70152015c0008fe2b006a01c7fffd;
mem[617] = 144'h0201ffd7000902280151fe7a004b0207ff21;
mem[618] = 144'h009b0225ffce02180265ffb4ffd702a202b8;
mem[619] = 144'h023200d705580029fe50fecbff4e00bd02a3;
mem[620] = 144'h012000b6ff6b0156ffb7ff0201d1febb017d;
mem[621] = 144'h01aafec6fe91ff2efe9c018901cffe790045;
mem[622] = 144'h01a600b6ff2bff4ffe97fe5dff07022700f2;
mem[623] = 144'hff4f000901ae00abff3a000f01a7ffce017c;
mem[624] = 144'hfe4b0023ff39fd75ffde012bff60fe7b0135;
mem[625] = 144'hff6aff130085febd0117ff7d011500adfe51;
mem[626] = 144'h008800d20122fde6006200270012fffb00f7;
mem[627] = 144'hfe8500100136ff57fefc0154ff60003dffb1;
mem[628] = 144'hff3afe73ffd50185012700bdffb3fdfc0167;
mem[629] = 144'hfecc013d0116ff0a0036014201a3ff11fdf3;
mem[630] = 144'h00d0ff320050007e01ba013b0000fee300af;
mem[631] = 144'hffd60010feb6ffdcfed201f001c8fedd0065;
mem[632] = 144'h01660157ff83017dff040089ff94ff9aff58;
mem[633] = 144'hfe3cfe590226013afe90fed201ebffad00cd;
mem[634] = 144'hfe26fe90fe1a00e2ff77ff8c0115fea901f8;
mem[635] = 144'h011b01e5fe16ff190176ffa8fe6e009a002f;
mem[636] = 144'h00cd0021feb1feb6fe4e003c018eff63fe47;
mem[637] = 144'hfe80fe6fff420195000ffe7c00d3fe2f00c5;
mem[638] = 144'hffbdfde00041fde7fef5ff240121fe4f0078;
mem[639] = 144'h0071ff020058fe4dff7d00ad00a7fdfcffbe;
mem[640] = 144'h017f02680556049e02f500e20236009001ba;
mem[641] = 144'hfef402e90340074e05190173025dfee6017a;
mem[642] = 144'hfff600b2ff8201db0268039eff9cfc40ff48;
mem[643] = 144'h01770439052e03b3023d000502f900effde0;
mem[644] = 144'hffcb019001f60173028501f3023500b4009b;
mem[645] = 144'hff8bfed20204fb34ff8502ebfcdf0057ff2a;
mem[646] = 144'h03d0054a03950090007c0206048ffcb90000;
mem[647] = 144'h017402c5fd41fdc1fbbb049902d6fe1ffe3a;
mem[648] = 144'hfecd0224027406c602670005020a022fff41;
mem[649] = 144'h027e031604df0308035802bc01d4fef2ff77;
mem[650] = 144'h02ea024904cd0311017fffb403750122ffbf;
mem[651] = 144'hfe27ffadfb4402b1ff0ffe16fdcbfc0dfe9f;
mem[652] = 144'hfde300caff3dffcdfeddfd7b00a8fe5bfea5;
mem[653] = 144'h00b50076ff07003f0059fe88ffd5ff4f0075;
mem[654] = 144'h000b015e033b05790610025a000a030900d4;
mem[655] = 144'h00dd032c048c065304b0009e01c401eeff84;
mem[656] = 144'hffdeff11fff3ff6ffeb5fdf800ec017c0000;
mem[657] = 144'hfe8ffe47ff2cfede014f018bff9d0179fe56;
mem[658] = 144'h01900030004601bf006cff94fe920085fe53;
mem[659] = 144'hff2600fe0119ff46fe6d0185fe3afdc0fddc;
mem[660] = 144'h009b0085ff25fe11fff8feb60112ffb3001a;
mem[661] = 144'hff47fe850138fde5ff4f0000013eff5bfefb;
mem[662] = 144'hfef5fe04ff7dfe9b006a010d0124ff25fe33;
mem[663] = 144'h002a0000007ffeeaffc4ff6f0034ffcf0086;
mem[664] = 144'h00aeff070031005afe75fed300ccffe000ee;
mem[665] = 144'hff32ff230081014a0050ffdbfdab0071012a;
mem[666] = 144'h00fffe2efe55ffa5023e022300fb0029fe7e;
mem[667] = 144'h010f00b70080ff6e00ba0060fdc8fecc00f8;
mem[668] = 144'hfe53fe65000dffd7fe880036fffdffdaffd0;
mem[669] = 144'h0063ffde012dff1d015cfe4bff14fe31ff52;
mem[670] = 144'h0014fe94ff44000f004e007d00ba011c006d;
mem[671] = 144'hfff8ff970118006dff63fe6701350139ff60;
mem[672] = 144'hff1e018afd9603950362ffe6fe92fea9fcab;
mem[673] = 144'hfd4bff72ff6503a902730254fe42fcd6fe71;
mem[674] = 144'h0338ff33fd05062c06c208630726017201e5;
mem[675] = 144'h0117fe3cfcf400760141011000edff1effca;
mem[676] = 144'h00edfd29fe140236039801bd0090ff6300de;
mem[677] = 144'h00a00094007c00af04b207b4068d01a7015b;
mem[678] = 144'h0052fb7ffb6302a2060e057ffe1d02b20174;
mem[679] = 144'h04ddfb15feda013108180ecb05a305f402a7;
mem[680] = 144'h002f01b5fd6003250390fff5fed8fd39fe3e;
mem[681] = 144'hfc86ff5afe7c02a004db003cfe1afefffe73;
mem[682] = 144'hfef5ffe7fd2b02b505db020202d1fe2dffa0;
mem[683] = 144'h070601860253ff39fe8a02be0727043403c2;
mem[684] = 144'hff58ff5a00e300a1ffc4feaffe38feb10052;
mem[685] = 144'hfeb6007f01ad006dff56ff2200b7009b00d4;
mem[686] = 144'h0129042dff4b01110000febefeebfe55fd10;
mem[687] = 144'h0116003aff17034a03760330002dfc91fe83;
mem[688] = 144'h025101b701c005240266fcd5fbbb000404ad;
mem[689] = 144'h02dc011800f7044101bffe4afc2202250477;
mem[690] = 144'hfc80fe4f046e05080329ff1a01130306020b;
mem[691] = 144'hffba0151039a02b9038afffff9ea03bc0319;
mem[692] = 144'h02e00080037803e80095fe34fbf0031a04d2;
mem[693] = 144'h0166fea001b5ff6f017f035ffdf2ff8f0116;
mem[694] = 144'h019507be06d6006f02ddfd0fffe20158ffe9;
mem[695] = 144'hf961050a033701ab041d04b202f8fdfbffdd;
mem[696] = 144'h01b60102037402d101d8ff04fbc601040358;
mem[697] = 144'h023c034401b7007e0155fdb2fc7201b20635;
mem[698] = 144'h02b4032202cf004c009aff16fd0c00ae02f3;
mem[699] = 144'hf979fa80ff0c02f701fd00e404850284ff75;
mem[700] = 144'hfe3800ef01550091ff72ff50ffed001fff31;
mem[701] = 144'hfe8501b9fe80009800bc014dff02018e01aa;
mem[702] = 144'h046f0108011b037902b7ff39fcf60225030c;
mem[703] = 144'h01bb01350201031700d4fe0bfe89001d03a9;
mem[704] = 144'h016c029c03de00d4fcadfdc1fbb102d105f4;
mem[705] = 144'h029803d00345fecdfcd6fffffc9901ee05a1;
mem[706] = 144'hfb9803450469fd700117fe75fd81051fff56;
mem[707] = 144'hff7601ea0221fe77fee001f4fe1efff803bb;
mem[708] = 144'h00d7008c0401004cfed0fecefe0101c7008b;
mem[709] = 144'hfc60000700a1ff35fd3ff949ff7efa46ffb8;
mem[710] = 144'hfc73055003b4ff0300520246fbd3fe63ff2c;
mem[711] = 144'hf7d6fe250009fd0e01e002ebfd6efda4fcbc;
mem[712] = 144'h015a02eb03f8ff78fdc8fed1febe006703ce;
mem[713] = 144'h010d039d04abff69ff1b000efc50023e06b0;
mem[714] = 144'hfd57015e03ffffae0033fe94fc62fde80287;
mem[715] = 144'hfa94f885fe60fd37ff47fbe5fdc90182fd4e;
mem[716] = 144'hfffcfe9000c501d60034fdaaff7a006d0169;
mem[717] = 144'hff0800c900edfe86fe6eff81019fff74fe36;
mem[718] = 144'h01c501d601e2ff92ffe7fe7ffdd3032b058b;
mem[719] = 144'hffea0182019bfde9ffc2ff1afc4a000204c4;
mem[720] = 144'hff46fc18feb2fe940220020f024b03680313;
mem[721] = 144'hfe45fc74feefffff0291ff6f00b403e403bd;
mem[722] = 144'hfd3a017a01ab00e2fd2affe6043c04c40084;
mem[723] = 144'hfad4ff18054b0294fe8c01c50476067d0111;
mem[724] = 144'hfe59ff36043d00dbffaeffc3049705ca03ae;
mem[725] = 144'h038f00c60116ffce051202e30052060401dc;
mem[726] = 144'hfe91062e0333feadfcf102a7064b0425ff6e;
mem[727] = 144'hff770557023a0041facfff6e086d00bb02e6;
mem[728] = 144'hfd84fd34029f02c4013e0180020201e2034e;
mem[729] = 144'h0100fd01021afc8f025e015c04e200fb0142;
mem[730] = 144'hff81ff7000dc0032ffe202a002bb065100dd;
mem[731] = 144'h0173089c02e502ccfde0030e055f01280288;
mem[732] = 144'hff7301310260ff800128fec301baffe20101;
mem[733] = 144'hffd900be0077ffe8fe80ff65ff2a00f1fe6a;
mem[734] = 144'hfedffdeefe980136016bff4eff7400c20262;
mem[735] = 144'hff1dfc190247ff73000c0246006f028c0225;
mem[736] = 144'h0066ffa7ff07ffa8fdc200da0164ffc9002a;
mem[737] = 144'h00530082ffa1feaf00e6fe260033fef500d8;
mem[738] = 144'hffda0160fe5dfe22016200e601beff5afe99;
mem[739] = 144'hfea5fdc300b4fea0ff6b0128008cffd2002a;
mem[740] = 144'hffa500ef00280154ffa1fecd0069000a000d;
mem[741] = 144'h003200bf00e6ff7f0108ffc300dbfe7eff09;
mem[742] = 144'hfe81fed8fe4affd2ff3ffdbe0075000c0158;
mem[743] = 144'hfee3ff39017e00cbff0dfe1afdfcfe6d000a;
mem[744] = 144'hff66ffc000c1fed5fed3ffd6fe200034fdc3;
mem[745] = 144'h007b009dff490054fe6f00c400da00ba00ea;
mem[746] = 144'h017500dffecbffacff5b0038fe8f00b300fb;
mem[747] = 144'h00d3fff3010bfe63fe9eff54ff50012f0143;
mem[748] = 144'h016600d0017e00030092fe33ffdefefb013b;
mem[749] = 144'h00600023ff47fed0011bff48fe35011f01ca;
mem[750] = 144'hffd5fffdfdc8ffa5fec5ff99ff58ffcd003d;
mem[751] = 144'hfeb3ff3efe83ff7200c3fe5e010dff24feb4;
mem[752] = 144'h01cf003d044d00df00ea00c200e4ff4cff88;
mem[753] = 144'h016c00ba02ef03140150ff9c012c00cafef6;
mem[754] = 144'hff0afeb9ff99fe42fae3ff84fbd5fb79ffec;
mem[755] = 144'h00a701740259002e0041feb00306fdddffe3;
mem[756] = 144'hff50017b00530005fd3701bd00effd76ff56;
mem[757] = 144'hfe7e0082ff5ffec301f5fd0bfedc024dfeb2;
mem[758] = 144'h00c9024e01cffde0fd5cff220327fe9efe4c;
mem[759] = 144'hfe1e025f0123fcb7fd52ff96fe7dfc41ffc4;
mem[760] = 144'h01d7016a015a0131ff7b0244021ffed3ff68;
mem[761] = 144'h028bff3e0325fd7e00fc00a0042d0082ff72;
mem[762] = 144'h022e0244012000e9fdc8fe9103d6fe18fdfc;
mem[763] = 144'hfad6fef4000102d6fe750313fc8afe5f0092;
mem[764] = 144'hff720043fec3fdeb0011fee3ffe501effde9;
mem[765] = 144'hfe9c006afe3ffe62019afeb700ba0124ff78;
mem[766] = 144'h02b400f404f603c305370073004a0280ff1d;
mem[767] = 144'h0138012802c8028400670106005ffeeaffe5;
mem[768] = 144'hffd7febd0064ff0c02a6ff300012fc0001f8;
mem[769] = 144'h025cfffdffea01830121ff8eff8dfe6d005e;
mem[770] = 144'hfe27feba058401480176fdf5fd2cf7d70280;
mem[771] = 144'h018dfe65010f013a0315ff07ff4cfdb001fc;
mem[772] = 144'hff76ff3f020600f00220fe4eff58fdb501f8;
mem[773] = 144'h0327fb11ff5102d3063b061f018bffc4000b;
mem[774] = 144'h01e405ba039f01ff0001fc2eff5c02090006;
mem[775] = 144'hffdd09ae0415025f009cfdecfefd009800b1;
mem[776] = 144'h0250fec300410278013a007c013fff3b01e5;
mem[777] = 144'hfec0fca10066005ffd7bffa400960136013b;
mem[778] = 144'h001dfdbb02930252fedffe6afde700bcff03;
mem[779] = 144'hfc1ef609fcfa032f00e103140107fcdeffcd;
mem[780] = 144'h002700000109003bfe1600ff00aa01c2ff2d;
mem[781] = 144'hff9b016600f5fe3d01970138ff61fe39012c;
mem[782] = 144'h0014023a03f3022effc2018500b100a3ffe8;
mem[783] = 144'h021aff4d0204ff26ffd6fedcfeffffc20047;
mem[784] = 144'h03cb03ad04430159ff140039fefe02530551;
mem[785] = 144'h039b03ad02b2ff850180ff9cfe6903a403d4;
mem[786] = 144'hfd6c003d0210fd5efe79fec0ffac0229ffc5;
mem[787] = 144'h013e034a05a800980102fe1f016604ab042b;
mem[788] = 144'h03c203d102fa012eff82ff44011901710282;
mem[789] = 144'hfeca0296040efee6fbeef96afee1ff320089;
mem[790] = 144'h01ea0902074bfdfefe7504bdffe3011a0253;
mem[791] = 144'hfd5e0319018bff5c01a00348034afd57fef3;
mem[792] = 144'h0454046f0124003000cbff47011b026404b8;
mem[793] = 144'h046406f80461002c01500154fd0c05930585;
mem[794] = 144'h0241042803d1ff1bffc00063004501a10498;
mem[795] = 144'hfad9fa5b00dbff34ff2bfb3501feff73feb2;
mem[796] = 144'hff7bffe60083ff2a01c5018200b800c50127;
mem[797] = 144'h01a900d20036006efe8bff0efe8d01b7ff43;
mem[798] = 144'h029202deffde028200a0000202d9056304c3;
mem[799] = 144'h030f03050380003001620159fe7104640398;
mem[800] = 144'hff0efe0200220046ffce0005ff29fe0d00b2;
mem[801] = 144'h00c501c4feb8006e00a30110ffcc0127ff17;
mem[802] = 144'hfd36ff4afdb5006eff10fefbfe3fffd8006f;
mem[803] = 144'h0029fdc7ff240112fe040011fe52fe3ffe0b;
mem[804] = 144'hfe87ff71fda900abfdc70028feb500c1fddf;
mem[805] = 144'hfee0ff09feb5ffcc0070010afe54fead008a;
mem[806] = 144'hfff1ff2fffacfea80064ff650085ff87ffbf;
mem[807] = 144'h00cffe47ff220087fd8e006ffeb3ffbaffcb;
mem[808] = 144'hfe46ffecfe82ffbfff5bff5f002eff020069;
mem[809] = 144'hfed5fec3fe8aff260120febcfe660151ffc2;
mem[810] = 144'hfd85fe52febf0064fdc5fda9015600edfe3d;
mem[811] = 144'h00a800c70029fe53fe5afef600650075fe03;
mem[812] = 144'h016dfec1ff82fff9018cfe7f01c0017f01a7;
mem[813] = 144'h016effe2ff8001590039ff180194ff2f00f0;
mem[814] = 144'hfdd3fdd7fe4cfdfaffc4ffe4ff70fe63fff9;
mem[815] = 144'hfeb8ffa90074fe3d00d6ff9eff23ffceff1b;
mem[816] = 144'h00e7ffe6001106e8020dfe25ff62fc3df90d;
mem[817] = 144'h0366ffdcfe4d05bd016afed7fdeffed5fa2b;
mem[818] = 144'h0386fd07fd6c05ad05a7041302abfea9032c;
mem[819] = 144'h04aa028cfae303eb02c302cafeb4fdde0108;
mem[820] = 144'h024a01c3fccb042e03440256fdd0fdab00ed;
mem[821] = 144'h05e10052009f01e3055e057f01ee02370016;
mem[822] = 144'h01c2fb8bfde1055305ec028c0080ff5c0252;
mem[823] = 144'h0174fef6fe70039d07540999053405e3029a;
mem[824] = 144'h0232029affb102d200bdffacfe88fc33fdfd;
mem[825] = 144'h0158ffefff52055c0110fd3cfe50fc22fa76;
mem[826] = 144'h00d1ffd0fd0b064c05bb008b00c4fd83fed1;
mem[827] = 144'h042d0155011301fa00c600e002e1ff1203d7;
mem[828] = 144'hfec701eb007001d7014f013fff4cfea2ff8e;
mem[829] = 144'hffe9feffff47fe31feb30176005c0112fe1f;
mem[830] = 144'h02f10158ff2001b800e3ff7affe9fd6afbc5;
mem[831] = 144'h00c70246fe8002b803bd01f1ff41ff56feae;
mem[832] = 144'hfdf1fe4bfb89feadff4900cb00a2febefb5e;
mem[833] = 144'hfecafec5fbdffd70fd9a00aa0264fdd3fd92;
mem[834] = 144'hff54fc39fae6ff9f0037fddb028b039b01f6;
mem[835] = 144'hfebdff9cfc6a0017ff95ffcb00f4fefc00a6;
mem[836] = 144'hfee9fd1bff4b007701c3ff7e01c3002500e4;
mem[837] = 144'h04c40311ffce0378055a04130743036cffff;
mem[838] = 144'hfe46fb45fd7b012500d9fec601c001a60329;
mem[839] = 144'hfd27fc3c00ab047d020dfc5cfb2202d20395;
mem[840] = 144'h00b9fdb7fd32fcfdfdbb0058ffe2ff02ff43;
mem[841] = 144'hfe29fd28fce2fe3dfe2eff6003d4fd15feb8;
mem[842] = 144'h00b4fb4ffc19ff4cffe8fe63003d0034fec1;
mem[843] = 144'hfd5d0756057a0000049807cd01910313028b;
mem[844] = 144'h009c00330078ff7ffe48fe7000ef01cd020e;
mem[845] = 144'hfef800c4feac00fbff41ffae01b201700083;
mem[846] = 144'hfdb9fd19fd52fdf0ff1a0010000cfce9fe6d;
mem[847] = 144'hffa1fef5fc78fee9fe55002d0202002affbe;
mem[848] = 144'h018301ad0191fcf901cd011c0058ff28fd67;
mem[849] = 144'h021d0312002eff4c000f036902ccfe19fb6d;
mem[850] = 144'h021efe5c02d1ff15fe70ff8bfff7fd890142;
mem[851] = 144'h039dffb8ff26fe9affa601d0ff3ffe5ffecf;
mem[852] = 144'h02db0020ffdefdc4fefb00c20182ff60fcaf;
mem[853] = 144'h01420047015fffa5fcc7fe7afe7aff7aff78;
mem[854] = 144'h0424fbf2ff54fef5ffee00b4fef2018a0164;
mem[855] = 144'h057e00c0fe82004dffcdfe2f0289056c0121;
mem[856] = 144'h012d00af00a1fe38008b01410299fd4aff10;
mem[857] = 144'hffd8fea001bbfff6fe150204001cfdcafb86;
mem[858] = 144'h02ea01acfe14ff96ff62ff4d034800c9fddf;
mem[859] = 144'h0223ff0dfff600700159012bfa1bfb5100c5;
mem[860] = 144'hff88005d0208fed6feb1017f003b001701c2;
mem[861] = 144'hff8d0169fe72000dfe4a018e019afe9c01c7;
mem[862] = 144'h008c00e402abfcf7feaf043201f8ff7bfc26;
mem[863] = 144'h0185001efff7004001b0027f00c8004aff05;
mem[864] = 144'h02700181012701d6026b05100259015c01ab;
mem[865] = 144'h01bb026f03a30296005b0222030201550137;
mem[866] = 144'h035f02dc033bfc0900c7fcdbfcecf937ff35;
mem[867] = 144'h045a0260040001af01e300220307fe960036;
mem[868] = 144'h0493028e014d00c0ff29005b038efeaafe13;
mem[869] = 144'hfce9ffb3014b0059feebfbbffcadffb20072;
mem[870] = 144'h043702ad022dfe96fc8a007002adfe55013f;
mem[871] = 144'h05ca057c0082ffb8fc12fcbdfc64ffa3fff1;
mem[872] = 144'h0199ffc603a502ad00c4028601dc01bb015f;
mem[873] = 144'hfe73010b00c60055feae00210283feca015a;
mem[874] = 144'h02f6011c011effa9fe24fef9ffcafeb1fca0;
mem[875] = 144'h0077fab7fd0dffbe03d5fd0af6f2f82afee8;
mem[876] = 144'h00da018501790262ff7a01a6ffcbff1501a7;
mem[877] = 144'hff6cff28feccfe66000cff7900fc004afeca;
mem[878] = 144'hff6c021102db016302d505ec047d03a202e6;
mem[879] = 144'h02f2016201e702b4fff601ce01aa030902d1;
mem[880] = 144'h02ba01460079039601fb04190142022204af;
mem[881] = 144'h044d0423016602f104bf028eff7a01e20272;
mem[882] = 144'h01c701b603e3fda700f4fc5bf5cefac700cf;
mem[883] = 144'h0521036c0163007400c2ff1a004c014e0054;
mem[884] = 144'h041e0434026dff9c020dfed8ff4c0186016a;
mem[885] = 144'hfddbff0d01befcbef91af912fa22fd94fec5;
mem[886] = 144'h040608810401fe6dff12fc98fb96feac012a;
mem[887] = 144'h03920510021cfe4efdf2fb4bf8c4faebfc66;
mem[888] = 144'h041202b1010801970189012b002e01f100d8;
mem[889] = 144'h016803820224fec800810115011f01d6049d;
mem[890] = 144'h01a3025803e0ff0b003dfec5fd1b00dc019f;
mem[891] = 144'hf9c7f432f8f40245016bf903f930fc80fc42;
mem[892] = 144'hfe390009018201ba000dfea4ffefff760166;
mem[893] = 144'h00d90060fff9004dfe0ffe69ff07009eff22;
mem[894] = 144'h015302ab020d03d7041803f400ee03ef03ee;
mem[895] = 144'h033b01d30045028103b102bf006304750256;
mem[896] = 144'hfdccfa5df851fd86fd100207fdd1fc52f969;
mem[897] = 144'hfca8fa6ff809fc4bfd3bffa7ffdbfc20fd2b;
mem[898] = 144'hfe66fa58fdb400c0007c021d05b105fb015d;
mem[899] = 144'hfcc3fa6bfb17fd8dffc100c4ff5f002601dd;
mem[900] = 144'hff34fbdafae6009701ecffce017f00ae0186;
mem[901] = 144'h04f7012bfc5701d5048c0564083200ee00b5;
mem[902] = 144'hfa99f90c008f01b502bc02680518060c01bf;
mem[903] = 144'h0069fe5902d7046d03fe01e606210b1c03ff;
mem[904] = 144'hfe49fc0ffa1afd18fefb023a0014fe23fd9d;
mem[905] = 144'h0041fb90fa6cff0dffa800690140fda0fbbd;
mem[906] = 144'hfe56fd52f9f100a9fffb0017ff9f00bffea5;
mem[907] = 144'h043103f006d2023301a7030b01230713031f;
mem[908] = 144'h004601390032fe2aff1000c3005a0069fffb;
mem[909] = 144'hfe2effd2019bfef601abfec101e200edff05;
mem[910] = 144'hfe11fd0ffa1cfdd8ffc000b0fd2cfa66f916;
mem[911] = 144'hfebefcdefbbefd24ffb60248003dfe07fd8a;
mem[912] = 144'hfe38ff13ff9b003c0043ff970028fecc0113;
mem[913] = 144'h00a3fe31fdf5fe67fef500d9fdecfefafe0e;
mem[914] = 144'hfe4e0050febd00a0fefcffd60058ff3bfe93;
mem[915] = 144'hfdc7fd730008fde0febeffc5003c00a3fdef;
mem[916] = 144'h00b6ffaefe17fe92ffc400ddfe94fdc6feb8;
mem[917] = 144'hfeb1fd7efe09fec400d8fdcdff9900cffe89;
mem[918] = 144'h0093fed0fd95011afd9bfef5003c0073ff06;
mem[919] = 144'hfd9bfffffe26fdedffb1fed0ff5dff8d0050;
mem[920] = 144'hff85ffc1fddd0069ffd0fd73fea9ff54fdea;
mem[921] = 144'hfed20077ff7d01150127fe780028fe2bfeee;
mem[922] = 144'hfe2dfdf8fee1005ffe4dfea100edff38fdeb;
mem[923] = 144'hfd7afee7010dff620113ff80fe920000ff65;
mem[924] = 144'h0108fe65010fffed01d50143feb9ffdb0124;
mem[925] = 144'h0038fe3301280127011101a4fedf00ea0028;
mem[926] = 144'hffdfff33ffac00310065fda8fea5feb2fda1;
mem[927] = 144'hffa501250018004f0046ff2c0068000efe04;
mem[928] = 144'hfd19ff43ff8dfc3ffe7002270042fe27fffc;
mem[929] = 144'hff7d001cfde7fca8ff9f019001b9002c0165;
mem[930] = 144'hfd64ff18fc90fff2010bff56fb8200e5ff3a;
mem[931] = 144'hfcaffc07fef3fba0fd8000780271018100c3;
mem[932] = 144'h0005fbf90042ff25fe3a0328ffd90178ffd6;
mem[933] = 144'h0213fd8e002f00de00eafd2b059a00e3ff53;
mem[934] = 144'hfae4fc2ffeddfc79fcbeff780175fdc4fd7d;
mem[935] = 144'hfb98fba7008cff16fda0f47ef837001dfd98;
mem[936] = 144'hffdbfef2ff4dfb55fd2f0160017bfeb0fffb;
mem[937] = 144'h0031ff1cfeddfdc50017040d0076ff0c0183;
mem[938] = 144'hfcd0fe3bffe1fcdafe1102f8016dfef3013b;
mem[939] = 144'hfea9014dff10ff77025c04b7fb6afff0fdca;
mem[940] = 144'h01ed00460270ff83fe01ffa6ffb800f7015c;
mem[941] = 144'h01adff3afed40118fee0fe7c00fc0158fe4a;
mem[942] = 144'hfeacff35fd66fb8afc90fedf01d3fe88ff82;
mem[943] = 144'hfe75fe4f0045fbf6009500f7009bfefe012a;
mem[944] = 144'hfda4005e0057ff9500430112fd8dfdc3fe03;
mem[945] = 144'hfef10034007fff3c00a2fd6dff7100e7ff25;
mem[946] = 144'hfdd9fe2b020dfef1fea2fdb6ff69ff8fffb6;
mem[947] = 144'hfe52007fff90fe23feda008f00a8fe93002d;
mem[948] = 144'hffbbfe13003200fffddbfea9ff39fe7efd97;
mem[949] = 144'hfda2ff220061fd85fdf400aaff03fe5ffef2;
mem[950] = 144'hfe93fedeffefff59005bfe0600bafdc5ff80;
mem[951] = 144'hffb7004900ffff0ffe5200e1fff3ffa9fea2;
mem[952] = 144'hfd90fe61ff1afee4ffb3ffc0fddafe690115;
mem[953] = 144'hfea90076fecf00f400490124feb40059002c;
mem[954] = 144'hff1500f5fdcf00f1ff08fd7c0054fdadfe80;
mem[955] = 144'h00ec00e00112fe800030ff3cffed00a90055;
mem[956] = 144'hffb9014cff1dfefbffd10040ffdd001f00eb;
mem[957] = 144'hff9301a1fe2500d1fe2affa901ab00c8fe82;
mem[958] = 144'h00f0ff530035fde6feb8000cfd8700d60120;
mem[959] = 144'h00c5fe13ff5afefafe10009800c9fdc7fefc;
mem[960] = 144'hfdcf01070125ffc30149fdc4fe0200f4003c;
mem[961] = 144'h0023010aff23011700e0ff6d0101ff2cfeb0;
mem[962] = 144'hfdd9fe4aff14fea40097fdecfe74fe49009b;
mem[963] = 144'h00e2009fff66fe400111fe11fdeffe78fe5c;
mem[964] = 144'hfdd2006d00f201760071fee80038fe85003b;
mem[965] = 144'hfdbfff9dff2b015a0078ff6500e30052fdff;
mem[966] = 144'h01530029fee3001801760024fe33002f0048;
mem[967] = 144'hfee2fe57fee7fe590137010c0077ff570153;
mem[968] = 144'h014c007efebfff5300580086ff94015cffcd;
mem[969] = 144'h01c8ff89ffb3fe1affc5ff41ff48ffdafe45;
mem[970] = 144'h01660017016f005bfe9d0084ff4efe4c00c1;
mem[971] = 144'h013501a7011500d00007fff5fe3e0195ffe5;
mem[972] = 144'h006ffe7cfefa018b0016005f00c00138ffe3;
mem[973] = 144'hff32fe6afe8f017dffa5ffd9fe66ff2cff49;
mem[974] = 144'hff59005d01190014fe2a008b00c7febcffc4;
mem[975] = 144'hffd4ff71007100eb00120116fedafdcafe62;
mem[976] = 144'hff46fe7ffd3fff48ff3efd61ff88ff96feea;
mem[977] = 144'hfd04fe92ffd30047ff4efe5b00b0ff7bff1f;
mem[978] = 144'h0070fe44fe15fdf10006feb200a5fe7afeb9;
mem[979] = 144'hfd2ffe16ff26ffb6fdf2007b006dfeaa0082;
mem[980] = 144'hfd25007cfffd0054fd4afe440060fddafeca;
mem[981] = 144'h0057ff1ffce9fdf50397fd0ffd6ffda4fdb2;
mem[982] = 144'hfe5bfdabff9e0065fdaefec0fe45fdc5ffd6;
mem[983] = 144'hfe18feeafdfffdd5002f00d8fecdff51fe29;
mem[984] = 144'hff88ffaa0176fe7dffddfe0afe6dfd55ffa4;
mem[985] = 144'hfd12ff64fe8100a7fcbdff7afdcefe54ff69;
mem[986] = 144'hfe79fce2ff68fedffff8fe4cfe5efe9a0168;
mem[987] = 144'h016dfce60041fe60fd39feac0029ff4cfd09;
mem[988] = 144'hff19ff7ffe37004f01da0022fe46fe900059;
mem[989] = 144'h00610030017f0093ffacff7bffb800000144;
mem[990] = 144'hfd94fcf1ff13fda6fff1fea4fda7ff10fd35;
mem[991] = 144'hff5efdbcfe6cfd1d0018fcd1fd15fd2000c0;
mem[992] = 144'h0311046b02cb030eff7cfc9f000a020d01ad;
mem[993] = 144'h049001e400af01dffee9fefcfd3201c30168;
mem[994] = 144'hfe1efe2705f0ff9101cefb47fd30fc6302cf;
mem[995] = 144'hffc9011c0366016d01ecfdaffd78ff280065;
mem[996] = 144'h013d019a02a301b3ffc2fe8dfeac00a9012e;
mem[997] = 144'hffaefef3029f01320253ffc0f976fe800156;
mem[998] = 144'h036306e60323fef90177fd61fe37ff230007;
mem[999] = 144'hfafc071f034eff8501b200bdff75fcf3fb88;
mem[1000] = 144'h0588042e01df00dcff24fe59fe6b01cc043e;
mem[1001] = 144'h02d80585022c03530170fc09fe1e047b02ad;
mem[1002] = 144'h040201a702f501920109fb0bfcab010b03b7;
mem[1003] = 144'hfdb7f510f974fdf5ff48fc970266fda3fef2;
mem[1004] = 144'h017cff6c013500660058ff360015005dff50;
mem[1005] = 144'hfe25fe4fffe00107007d0100003bff3001a6;
mem[1006] = 144'h03800150035703a5005000700258027f0442;
mem[1007] = 144'h04c8042d01a00348021ffe7cffda017a01d0;
mem[1008] = 144'hffbafdff015403130289ff63ff18fd070354;
mem[1009] = 144'h0009008901c60190ffe4ff53fd3a000c01ed;
mem[1010] = 144'h03d70203047e041d0672071304e407550014;
mem[1011] = 144'h010afe42012500b501b901b9fe3000aa038e;
mem[1012] = 144'hfe80fcff022d035d02770351ff500146044c;
mem[1013] = 144'h04fe001d010b025a018f06d2061701b600b1;
mem[1014] = 144'h0093fc5501d5028d0668033202bd0566031e;
mem[1015] = 144'h038901f3020404b505430b5e06cf075d00e1;
mem[1016] = 144'hfec1fd600050ff95026f02610015fe1c0139;
mem[1017] = 144'hfe68000001bc01a3011401e0fdec003c02ad;
mem[1018] = 144'hfe86fd6201d70398041400d2fecfff140331;
mem[1019] = 144'h057e02bf04d003510106ffc705e30cfb0395;
mem[1020] = 144'hfe77014effa2ff6901ed0031fe71ffea0139;
mem[1021] = 144'h01430097ff7500e1fee900d2fe210183ffd5;
mem[1022] = 144'h021dffb5ff2b00a70027feeeffa4fbebffcf;
mem[1023] = 144'hfe3ffebc01fc021cffc101a2004bfefa033c;
end

always @ (posedge clk) begin
	q_a <= mem[addr_a];
end

always @ (posedge clk) begin
	q_b <= mem[addr_b];
end

endmodule