`timescale 1ns/1ns

module wt_fc1_mem1 #(parameter ADDR_WIDTH = 11, DATA_WIDTH = 144, DEPTH = 1024) (
input wire clk,
input wire [ADDR_WIDTH-1:0] addr_a, 
input wire [ADDR_WIDTH-1:0] addr_b, 
output reg [DATA_WIDTH-1:0] q_a,
output reg [DATA_WIDTH-1:0] q_b
);

reg [DATA_WIDTH-1:0] mem [0:DEPTH-1];

initial begin
mem[0] = 144'h04a40433fa38fea4fec6fca6fee003e30796;
mem[1] = 144'h04c3025ffb8a0014fcccfbb2027102b5064f;
mem[2] = 144'hfcfdf597ecf9002900bf030c0713046b005c;
mem[3] = 144'h019701cffae9ff9eff82fdfb010804c40309;
mem[4] = 144'h046e027cff4c02d80097fd8000650454029f;
mem[5] = 144'hffb004bd05a8fc280406f58ffcc200af054b;
mem[6] = 144'hff8cfde7fa110042ff0b010efeaefdf6fe2f;
mem[7] = 144'hf63cf67cfa7a00060073059d0215fa33f7e2;
mem[8] = 144'h039100f4fba0ff24fefdfbcbffa6052002bc;
mem[9] = 144'h038502fefc1a008aff59f8c9fe97035308f3;
mem[10] = 144'hffae0222fda1021d0014fe47ff1404590582;
mem[11] = 144'hffc2ff00ff2400fdfc01fe5106d90d91046f;
mem[12] = 144'h0042fcfdfd7702370208fe4afe07fe19fd32;
mem[13] = 144'hff3cfe8ffe89fecc0016ff83ffe001aa000e;
mem[14] = 144'h021afecafc7a040eff92fb12013904b5042d;
mem[15] = 144'h037d0313fd1bff49ffe5fdbd0068023d0483;
mem[16] = 144'hfe4c007600d100cbfe0bfe12febcffccff1c;
mem[17] = 144'hfee0ff54feabfe8c007ffdee007cff4aff01;
mem[18] = 144'h0178fe27ffa50071fe500216ff69016afe9b;
mem[19] = 144'h010bfdf0fe58fdc90061005dfe5cffdffede;
mem[20] = 144'hffcd00befe4400b90148008aff68017a00da;
mem[21] = 144'h021600910083fe74ff40fdfa00f5fdd7fef5;
mem[22] = 144'h009dfe4801b6fdc100a9fe140020ff77fdff;
mem[23] = 144'h00c3ff86003dfef5fe62fe8e008dffdc0048;
mem[24] = 144'h0052fe26ff6b01720006fffd007dfddbff09;
mem[25] = 144'h014e012d0034fe8fffbeffbe010f016bff48;
mem[26] = 144'h0147fe75017dfdfa0065000bffff01580214;
mem[27] = 144'hffc7fef801e2fed9fe380055017702390068;
mem[28] = 144'h01d0001aff9a019dff55ff07fe3a004bfee0;
mem[29] = 144'hff96fe58febffe2ffeed018e002eff95ff64;
mem[30] = 144'hfe96fe11016affa2fffe005c00d1ffcd00ac;
mem[31] = 144'hffb1ff8effb7fe2700d2002f00ae00e200d5;
mem[32] = 144'hffd70042ffed0047ffbeff88ffe0ff65014a;
mem[33] = 144'hff13fdd4ff66fdd100600175fee3ffff00c7;
mem[34] = 144'hff1fffe801310104ffe1feb1000300d7ff71;
mem[35] = 144'hff84007dfeabfe0300a3ff19fe6bffc6fe95;
mem[36] = 144'hfebf0184ffcf00c300c0fff00085ff2afdc3;
mem[37] = 144'hffd60014fe2c0021fed90037fed2ff41ff09;
mem[38] = 144'hfffd0026001fff2eff4cff8b002500150189;
mem[39] = 144'hfe5c00f8ff990096ffcffebefe1fff29005d;
mem[40] = 144'h00c4ff65fdffff6e003aff3b009d013bfe10;
mem[41] = 144'h0037ff80fef2014a007efe79fe5801db004d;
mem[42] = 144'hffff0111ff65ffe4febefed600ebfffc00c6;
mem[43] = 144'h01da01b3fe5d00d60121ffab006eff30fffd;
mem[44] = 144'hfef3016e00930166fe690057002a017c0029;
mem[45] = 144'h012b0038ff8fffe000a3ff18013300b3004b;
mem[46] = 144'hffa600590026fe4afe710015ffdffefcff0a;
mem[47] = 144'hffe4fe81fe5fffddffe600bf0040fddc00c2;
mem[48] = 144'h008b001bff0cfe9ffe7b0032fe12fdcafddd;
mem[49] = 144'h00b4ff04010100410096fe91fdceffbafe06;
mem[50] = 144'hfde5fff5fff1fff6016900e7fe87fe6c0092;
mem[51] = 144'hfd58fe73fe58ff8afe1bff49ff40fe3e00a2;
mem[52] = 144'hfe1fffb9fdbc00b4ff82ff66ffdf0109fdce;
mem[53] = 144'h01c60110ff18fed6ff4bffb900a80004ff44;
mem[54] = 144'hffa2ffd600f6ff52ffc7ff9cfe740037ffe7;
mem[55] = 144'h0115fec8fe98fdfdff6700070075008affbd;
mem[56] = 144'hfe60fecffd5dfe58feb5fef1fe3ffed100d9;
mem[57] = 144'hfeb6fd9c004efd62004efec4000eff52fff1;
mem[58] = 144'hfdfffdcdff3dfdc8ff7dff01ffe4fddb0078;
mem[59] = 144'hff6bfe7fff440107fedefe4bfee5fed3fea7;
mem[60] = 144'h0060ff440088010801250145fe3b0118fe82;
mem[61] = 144'h00e3002dfeb80154fee3fe830004012f011d;
mem[62] = 144'h0038ff8f002700e9fd6500b700bbfde3feef;
mem[63] = 144'hfda600c0febe00eb0042fdfbfda3feb4ffe7;
mem[64] = 144'h01a7036f037d05cd034a019cfe240207047c;
mem[65] = 144'h00c002450318022803ae0325ff37042f041c;
mem[66] = 144'hff57ffeffec4043e01d4faddff3307a302ed;
mem[67] = 144'h019004b004d402210548019bfdc8ff55ffea;
mem[68] = 144'h0192012d023b036102fe02f1fcc401e500c0;
mem[69] = 144'hfc1504f4021f004900300780fe1e046c003f;
mem[70] = 144'hff3403380018037400c0fc4efc83fa5cfd02;
mem[71] = 144'hf70ff6bdfa380400fd75f5fffc81f9d5fcde;
mem[72] = 144'h001c040f042b0270058d0242003701120221;
mem[73] = 144'h028402cc042f00a504780568fe13022a01f4;
mem[74] = 144'h018d03d90322017004d20310fe18017501a2;
mem[75] = 144'h06320ba302660351021bfa9d089311450399;
mem[76] = 144'hfe99ff67fe21fe2cfdc3ff88ff86fd9dfd50;
mem[77] = 144'hfe5bffecfe400070016ffe8a01b6013a0022;
mem[78] = 144'h004c00340273fde2026d034a00b6031e0305;
mem[79] = 144'hff2e01df02e203af05bf0341fe4a03d40468;
mem[80] = 144'h000f01b40033febbfde000860032fea6fec6;
mem[81] = 144'hff8bff59ff0901e10116002cff9dfe48ff5d;
mem[82] = 144'h00a6012cfffe017401bbfff6ff9efe5afedb;
mem[83] = 144'h00b600cf0118005cff090160009dff29fecd;
mem[84] = 144'h012000ad0136016ffdc8ff2b003e007b00d2;
mem[85] = 144'hfed3001a013b0086fe25015aff76ff5eff52;
mem[86] = 144'hfe9d007e016d004400b0fec20173fe41fead;
mem[87] = 144'hfe7c0150fdf9ff43ffebfdce006a011afded;
mem[88] = 144'hfeb8015100c400ab00e60033ff7bfe6cff61;
mem[89] = 144'h002cfe7cffcdfef00034fe77011cfebcffac;
mem[90] = 144'hff75fea201750196fe370135005efdde01eb;
mem[91] = 144'hffd0ff32014a001ffdf00134ffca00ccfecc;
mem[92] = 144'h01b60034fe70002aff59015efedfff8f00b1;
mem[93] = 144'hffb50121ffb3012000cbfe66ffd7015301ab;
mem[94] = 144'h006affe0ff010007014e00f2feacfe680129;
mem[95] = 144'h001afebeffdbff500001fe57fed5fdd8fed6;
mem[96] = 144'hfe0100e905f400ad016dffdafa2afbf502a7;
mem[97] = 144'hfcbc012902dd0235011a01d2fc3dfc010187;
mem[98] = 144'hfbe200ba0a360075ffd1fec0fbfffe820513;
mem[99] = 144'hfc88fe60043c020aff83027cfb32fc5d014f;
mem[100] = 144'hfcbafef50489ffcf01320416fbedfdaa0170;
mem[101] = 144'hfaabfa6dfff00065fe840853047afbdfff83;
mem[102] = 144'hfb1400df0741ff8102380011feb700f500d2;
mem[103] = 144'h005f03930321ffc5ffacfbb3046a036a004d;
mem[104] = 144'hfe69010902f300cc00a80240fa0bfedd0150;
mem[105] = 144'hfdd4011305e1fd8effd902fbfa85fed0011c;
mem[106] = 144'hfdddfc4501bafdf2029902d3fea4fd8c0116;
mem[107] = 144'hf9e1f902fbeb01090186fe83fccefce201f4;
mem[108] = 144'h01a3031f0149005e011effa30044002500eb;
mem[109] = 144'hfed80017018afe4cff6b009e015bff10ffb2;
mem[110] = 144'h02ed01d301f1ff110177011bfcd6fda802ce;
mem[111] = 144'hff7300200325014801ff012dfcc1fd7e024f;
mem[112] = 144'hfea0ff60fe44fe1d0007ff2ffee3fdf9ff5a;
mem[113] = 144'h0136fde6ffadfe20fed2013f00a6fe2e017b;
mem[114] = 144'h0077020c00db0115011ffdd201c1005aff1a;
mem[115] = 144'hfdde0030ff00fef5004100a40073fe9a0069;
mem[116] = 144'hfe24fe10ff38006c0049fe3c0077fe41feef;
mem[117] = 144'hff3500c60175014bff02ff9efed9015ffeb8;
mem[118] = 144'hfded02180102008c00c50124ff12fe15fe1a;
mem[119] = 144'hfe47ffd1ffc601360165002dff11ff3aff57;
mem[120] = 144'h0046fdcaff38ffcd0113fe6efef1fde9ff39;
mem[121] = 144'hff67fecc0133ff61feaa018f01380184fe9f;
mem[122] = 144'hffc5006800c100dffee6fdf500b700d6ffb6;
mem[123] = 144'hff67fff600ddffd70059ff6f0238fe27fe39;
mem[124] = 144'h0074013501810194009efe8efff8fe45fee4;
mem[125] = 144'h013dff40fed6fe71ff56006b001c0031ff9c;
mem[126] = 144'hfe43ffa6feedfdda010e012c017c0065ff42;
mem[127] = 144'hff970173ff05fe1eff44ff98016a0004ffd8;
mem[128] = 144'hfe33fe140113023f04ae03d805530408006c;
mem[129] = 144'hfe4c01fc0453034a04b50151024501c600bf;
mem[130] = 144'h04a90c0f07e00155fe9600ecff4dfd00ff82;
mem[131] = 144'hff3704be04af0231047c01e803ca008f00f0;
mem[132] = 144'h020403110366029f02bd0303018801ac014f;
mem[133] = 144'hfd24ffd00168ff3eff8003e6f65c018500a7;
mem[134] = 144'h0374ffc7018e0037ff08fdf4007cff270312;
mem[135] = 144'h07bc039201ccfe81fc56fb3cfedb014e01ad;
mem[136] = 144'hfe59004801960451025401d602b201c20049;
mem[137] = 144'hfe7b00cd02c704bb03ab01fcff7902a6fc9b;
mem[138] = 144'h0241013d01370347041e015700a902da0133;
mem[139] = 144'h05fa0b12ff4b02d70152ff48ff87f773fb40;
mem[140] = 144'h0038ff52ff69fd42fdad0273028cff44ff46;
mem[141] = 144'hffd500a5ffb0ffddfe5bfef6000d01130136;
mem[142] = 144'hfc8c01a505bc0271011c033304a001ae0022;
mem[143] = 144'hfe9101ac00600231025a0409030d018101f4;
mem[144] = 144'h04cb06c0038bfd4cfc93fd97ff5603f80155;
mem[145] = 144'h069a060a02e9fd85fe8dfc5d011f03a60092;
mem[146] = 144'h0139fb4ffa78ffa4007002c4ff6aff7f01a8;
mem[147] = 144'h049804d60352ff2afe4bff3cff98fcc2fa2d;
mem[148] = 144'h06c703b303abfeeffe9efe95fd45ff5dfe0f;
mem[149] = 144'h007e02cb02ccfe0bf794f92d001e00c9ff58;
mem[150] = 144'h07e403900099fe990181ff97fd2efdfefd49;
mem[151] = 144'hfce8fa63fcee0062042d05c6f99dfc3efd16;
mem[152] = 144'h04c1038c0276ff35fd15fe8b022f00acfed8;
mem[153] = 144'h089704ae0280ff66fe1dfda8febc01d5ff08;
mem[154] = 144'h051a044e0471fddafd0afe67fe02fefefbae;
mem[155] = 144'hf6cff8ea037cff79fc4501d60293029902b3;
mem[156] = 144'hfdd7005a002e0105ff140106fda40074fe6f;
mem[157] = 144'hfeef0078feae000c006c00a2013ffed9fe4c;
mem[158] = 144'h02c20517026a036d00adfde1049a031a01b8;
mem[159] = 144'h064805890312fea8fd84fc3201330095fee3;
mem[160] = 144'h00d1ff55ff3100ff01d90135fe9fffd1fbf7;
mem[161] = 144'hff69ff4b017302b30362ff86ff0f01fcfa43;
mem[162] = 144'hfd8efed4009b055006c2f8f8017afd37f936;
mem[163] = 144'h028f022b012700dd029b0000fc3f0401fd45;
mem[164] = 144'hff94ffb8fedefede014bff70fd900337ffad;
mem[165] = 144'hf95aff2cfcaa03aa02e90974fab805a1ff33;
mem[166] = 144'h010a020601c702d3015dfbac036c028f01c0;
mem[167] = 144'hffb902df007d0450035af9f104f5017e030b;
mem[168] = 144'hff820169002601a5043c002e00af031bfdab;
mem[169] = 144'h01de01bcff79002703100013fd3b04e1fb22;
mem[170] = 144'hfe6c018dfe86005003ac043afe6b027e0049;
mem[171] = 144'hf8a1f410fede00e90317fb1b0850f5c701b5;
mem[172] = 144'h02d700c301fbfeffff1400ff017a02e7ff46;
mem[173] = 144'hfe9fff71feab00edff1e009600000077ff73;
mem[174] = 144'h034d022700edfc7b014a02cdfca20011fb8b;
mem[175] = 144'h009bfff1013affdf03dd024ffcbc039bfe28;
mem[176] = 144'hfeb0fe7801c80219fe740099fea6ff6bffb0;
mem[177] = 144'hfef8fdd3021dfec8fffa00f9fdd1ff2c0174;
mem[178] = 144'hff4f000dfe7501550028fe6b023dff22005a;
mem[179] = 144'hfdc60087feccfec5012bfee4013301180044;
mem[180] = 144'hfdf9ff37fe2effa3fff5ffacfe3ffdcdff49;
mem[181] = 144'hfec2ff5efdda00ff0143fff6010affb200c6;
mem[182] = 144'hff5901bc00e4003efdcdfec3008f0142ff55;
mem[183] = 144'h016b003e0065fe14fe53ffd6fe660091ff00;
mem[184] = 144'h0109fe1afed90042000900f700c8ffcb0012;
mem[185] = 144'h009301510236ff9e007f00aaff9b0102ffed;
mem[186] = 144'h008dfeb00127016800edff65fe7c0153ffbe;
mem[187] = 144'hfeb500ed006bfe91fe680146fec4fe9e005c;
mem[188] = 144'hff3001b5ff87ffbbfe73fecd00140080005d;
mem[189] = 144'h01c000f7ff77ffedffc501940124fe23ff49;
mem[190] = 144'hfe04ff33fe8fffe6fe4d0069fdda00e9ff93;
mem[191] = 144'h0075010d0089fdd4fe88ff67fee3ffce01ee;
mem[192] = 144'hfeccff6f014000f101b1ffecff8a028d02c6;
mem[193] = 144'hfcadff170185ff0f011c01e9ff7a01b7021e;
mem[194] = 144'hff670641fd6e0097ffc7fdcd024302b7048b;
mem[195] = 144'hfbbd00c90030017cffb6ff1b00f30182023a;
mem[196] = 144'hfd6d01e3fea0fea6012301bc01f301d100e0;
mem[197] = 144'h01b301160103fc36fb09027dfacd0229ffef;
mem[198] = 144'hfeb1ff83fc1bfef20005010200c0fed800b4;
mem[199] = 144'h005800c5fa63feb40009fb43feb7008501b9;
mem[200] = 144'hfce9fe9cffb7fe0802c401010255fef800ba;
mem[201] = 144'hfb48fe92fefcfefd01bb0340ffe7fef800d8;
mem[202] = 144'hfd00ffd4023afe44016900e4007b029f0268;
mem[203] = 144'h0b5a114c03b4fe24ff8cfa120347039cfe12;
mem[204] = 144'hfdfd0040fe690176fda8fe2d013e0020ff39;
mem[205] = 144'hfe76012bff00013efec8ff48fe7dffeb004a;
mem[206] = 144'hfc02fdeb023702150211ffd2ff550058ffc6;
mem[207] = 144'hfe76ff870122003200bb01feff18008c0132;
mem[208] = 144'h025f0069fff500c5ff79ffa0024103b8fbf1;
mem[209] = 144'h03a5ff58fe9e033efeb3002a049100a9ffb8;
mem[210] = 144'h020602ebfc2802df00e6018f024f02a0fe45;
mem[211] = 144'h02320216feb601250317ff2302e1ff35ff03;
mem[212] = 144'h013602eaffac020e021fffb4031402c6febc;
mem[213] = 144'h09c2051000c1002102e800d10263037400d5;
mem[214] = 144'h02560000fb3d01450070fde3ff91fe58ff05;
mem[215] = 144'h01a5fda1fb8c009d006d03080063fdcb0109;
mem[216] = 144'h01d10112fe54015eff46fe1603c500eefc68;
mem[217] = 144'h02950091fe44017801b8fb6f02ac00d1fc7d;
mem[218] = 144'h03ba034fffc7026b0239ffbd022d016dff52;
mem[219] = 144'h086e101b0562000c005c02470b060cc80370;
mem[220] = 144'h006300b6ff25005600c5fdccff7b0174fdbc;
mem[221] = 144'hfe2eff83012d017101a6ffe001ddfef400db;
mem[222] = 144'h00dcfde9020d017a0076028401b1029dfe76;
mem[223] = 144'h038800bbfe070021fedd0030021802afff0f;
mem[224] = 144'h076c055903f1fdf0fda7fe3100cd02aa03f6;
mem[225] = 144'h048d065102e7fea8fd0ffd1bff98042003c7;
mem[226] = 144'hf978f629fa65fd7ffd9afd7dffeb02d5fae9;
mem[227] = 144'h047d03e10403ffaaff29fd20ff4002f1fd02;
mem[228] = 144'h046c033f0339fe06fe17fcfe0000038ffc16;
mem[229] = 144'hf4acfede02df00d4fc0bfa83fb71007701fd;
mem[230] = 144'h00ba0434035efe22fb59ffb3fec3fea4f969;
mem[231] = 144'hf990f85efeb8ffacfcd0027b009bfa21f8f8;
mem[232] = 144'h04b103e70234ff4a0000fdf1fe5c026800e0;
mem[233] = 144'h05ab04d1021dff56fecefc15fdcc01ebff16;
mem[234] = 144'h04a305dc0344fd1efe10fd96fd00025dfc69;
mem[235] = 144'hf113f25cfcd4fe7efd22fa03ffbb012bfe3d;
mem[236] = 144'h02b6fe0dfedd0180ffafffacffc9ff50fdca;
mem[237] = 144'h0073fe820116feadfee7fe7cff72fe6f0079;
mem[238] = 144'h0774055f00830084ffd1000202230283058d;
mem[239] = 144'h0417064602b0ff95fd33fee5011801f80176;
mem[240] = 144'hfec4fea803c7056d050503bb00140003025d;
mem[241] = 144'hfdc5ff3a026d0334051a038bfe93fc1bff85;
mem[242] = 144'h0180022d06f607aa020e0071fa52fc5efe28;
mem[243] = 144'hfe70005d020102d102d106efffb4ffc503ea;
mem[244] = 144'hff47fed3013f03d1058c0490ff9a001503a4;
mem[245] = 144'h00c1febefd76040709430b24062dfdf3fea2;
mem[246] = 144'hfe8502ea04a0058e00ddffaf01050313043f;
mem[247] = 144'h02af04cf052202e3ffdff9bbfefe03a9010c;
mem[248] = 144'hfe78ffd1018b047d05410665fccd00090191;
mem[249] = 144'hfcba0136030102d603f103cd007200c10398;
mem[250] = 144'hff4efe00ff8b05b3036f049bffc4fdb403c4;
mem[251] = 144'h037ef57efb0d0505067b087ffddaf9d40428;
mem[252] = 144'hffee0339fedafe21016502e0ffdffedafffd;
mem[253] = 144'h013301dbffae0022fe6d013801b90186016e;
mem[254] = 144'hff80012d02c5fdf5fdf30431004ffc670029;
mem[255] = 144'h009f014000cb03fc0446053afc8f00050200;
mem[256] = 144'hfed7fd4c026bfdbf00b904870302fd3afece;
mem[257] = 144'h00d5ff3101c4fffd00fa049d040bfd2bff50;
mem[258] = 144'h018b02370b24ff04fe3e05a2fd92f922fa04;
mem[259] = 144'h0041fe220197ff4ffd7303f00235fe770128;
mem[260] = 144'h0010fe4e001a0012001c04ea0415ff66fe43;
mem[261] = 144'hfc09fc0afaba02abff16fd7ffeb5fc2bfb7b;
mem[262] = 144'hfd1c00bf03f9fd47fffa064b05a4027d0282;
mem[263] = 144'h037b0a740450fec5fe0804f3006f05350397;
mem[264] = 144'h005dfe58014dfe0aff1a02b50318fcbafe12;
mem[265] = 144'hfc1afca7ff91fe70023703a2012ffdc7fb82;
mem[266] = 144'hfdf2fe8000b3fccffd9004a0057eff30fdb0;
mem[267] = 144'hf944f435fa180208009e042fef31e752f9cc;
mem[268] = 144'hfe100138ffaf00bdff89007e01b80132014c;
mem[269] = 144'h0047ff7300860159018f016700a4fe210189;
mem[270] = 144'h00c502bd03f0019cfee000d5005afec4ff79;
mem[271] = 144'h0047fd3dfeb0fe0afe90030600c7fccffc8c;
mem[272] = 144'hfc2afed9ff8a006703abfe85f9b1fe6e0212;
mem[273] = 144'hff03008dff7701fd0278003afa35fb1800c4;
mem[274] = 144'hfce7fbcd0958037e003dfc81fdfbfd8cfdca;
mem[275] = 144'hff6dfc780316ffdb00dafe78f9fd00af0365;
mem[276] = 144'hfcc8fe38ff8dff52022d01ecfb91001703b6;
mem[277] = 144'hf710f988fcbd0197058e072efec8fb96ff26;
mem[278] = 144'hfae602a3076b019c008dfd08008f07c501d3;
mem[279] = 144'h0185078508860368008ffd6206b10519ffdb;
mem[280] = 144'hfd23fd0101c300e5038c000dfbe3fcb30305;
mem[281] = 144'hfbbd00c50268ffbf00c3ff2ef97400b700d7;
mem[282] = 144'hfc85fbce0197fef40055011afc6affbf01a6;
mem[283] = 144'hf5f9eb86f9b5044b0254fd4bfcdef4b5fe72;
mem[284] = 144'h001f022801250084005d01ebfe16028c010f;
mem[285] = 144'h00aa002a00b40066ff6100410139ff6600d3;
mem[286] = 144'h048700d30109feb7014d0148fa55fd5200c8;
mem[287] = 144'hfd03feb9014f00a8027f0064fcaffcfe0373;
mem[288] = 144'h0118039a05e2ff060260049f01d70196ff07;
mem[289] = 144'hfee90064057c000b023a05b602deffa9fc69;
mem[290] = 144'hff9201270d820202015002c400260032fc17;
mem[291] = 144'hfdc002c9059b00a3006e060b07070222ff1a;
mem[292] = 144'h00dd008a01f8006702a504f703940017fcee;
mem[293] = 144'hfb47ff06fe5601e501d3014001a20285fc66;
mem[294] = 144'hffe3021905ccff81ff7005f90454fe5bfdc6;
mem[295] = 144'hfcd7fe0303c00078fbb8fcd8fffbfedf003b;
mem[296] = 144'hfeb0038b03ac01ab00b405ac03bfff5cfead;
mem[297] = 144'hff7c0119048cff8402fd071002a1fe76fc28;
mem[298] = 144'hfe5e0293024600860194056506edffd5fabb;
mem[299] = 144'hff48041efda602120335022af39cf699f95e;
mem[300] = 144'hffa7004c0089ff010141034cffc0028b0340;
mem[301] = 144'h004bff52018900e4008aff2ffeccfe3efe3e;
mem[302] = 144'hffbe01510433ff0fffed025201c100f10155;
mem[303] = 144'h003702060454002202940622040e015eff54;
mem[304] = 144'h0077fec9fd82feb9fdb2ffab00bcfe6efdf8;
mem[305] = 144'hfee2013cff740161ffe4ffefffa1ff4afda4;
mem[306] = 144'h0016006dfe46ff0cfe8efe90fee0ff23fe81;
mem[307] = 144'hfddbfe68ffcfffab00d60036feb6fe15fdcb;
mem[308] = 144'hfdedfeb7fec20128feb7fdb00051fec30118;
mem[309] = 144'hfe7bfedaff75ff9d01c200bdff030029008b;
mem[310] = 144'hff0effeffe0cffd400ecfe1400120107fe05;
mem[311] = 144'hff8e0146fde2fec401290136ff5400f000ae;
mem[312] = 144'hfe7effe2fdd4fe20fdcafefeff0ffe50fdc4;
mem[313] = 144'hfff0fef5fdeafe25fe34ff7e009cff72fdd5;
mem[314] = 144'h0050ffa3fddbfee2fd9cffc4ff69ff3dfde4;
mem[315] = 144'hfe210110fe9a0105ff7effea009ffeba0113;
mem[316] = 144'hfe4cfe6d01c3ff2bffd0fe3300860000ff5c;
mem[317] = 144'h00d0ffb1004b01bcffeafe9b005afefb017d;
mem[318] = 144'hfe63ff97fe34fffa011e0088ffcafde8fee0;
mem[319] = 144'h014800cffe03fdf0fe570048ff32fe4200aa;
mem[320] = 144'h02fe0009fe27038f0187ffd7046c0255010f;
mem[321] = 144'hffff009cfe7102e402b800ed031104330013;
mem[322] = 144'h04da02a5f82e042306e30429ff910140ff65;
mem[323] = 144'h01f10281fddf033100e203c4040d01d10053;
mem[324] = 144'h04430014fffb00ea040c0447021d01600090;
mem[325] = 144'h0ac607000099ffe90864041803ac05a7027f;
mem[326] = 144'h01b6002ffd8b04e1047201dffedf0102ff95;
mem[327] = 144'h0012fd1efcb204f003e6020bfe08febf00b9;
mem[328] = 144'hffc80127fd6a02ca02d30098042a02360165;
mem[329] = 144'h009901ecfee40445029400a7017402ac042d;
mem[330] = 144'h028a01a2fbf7050d035a031f027effea03c6;
mem[331] = 144'h12420c0d04e7016f014d04d509f4077906a1;
mem[332] = 144'hfd70fe94fe2aff1502d4fe69ff4c0032007c;
mem[333] = 144'hff00ff42013d01600173ff12ff44006c00a5;
mem[334] = 144'hfcc6ffa4fefcfbd6fce70159011e02dffd9e;
mem[335] = 144'h01e30094fd3a03e8030e01c2009500ff0058;
mem[336] = 144'hfbbafbcafffe02e1017002730308fe82fecb;
mem[337] = 144'hfc9aff0b01df01a602ab03200159ffb6fd23;
mem[338] = 144'h033a0bc10cb2018affe9fd11fef5ff4e00ac;
mem[339] = 144'hfe7501e202b203dd03e80437014801e801b5;
mem[340] = 144'hfccaff9900de036e03b703fb0157012801ee;
mem[341] = 144'h0386ff4efce100da00d508a5fa9702f4fe21;
mem[342] = 144'hff56fe6c026d0116014400290413009a04cc;
mem[343] = 144'h064106f80256ff7a0091f9b4017f07f205bf;
mem[344] = 144'hfb39ff8101f5036b03100503038c00f5fe4d;
mem[345] = 144'hf9e2fc67fec9037e043a075e02c10080fc44;
mem[346] = 144'hfc7b00a6002e01160137045e040a0299fe06;
mem[347] = 144'h09ad0be9ff63010005b2ff99ff28f486fa39;
mem[348] = 144'hfeaf02480188ff7aff5302ca002600330132;
mem[349] = 144'h00f0fe93fef2fe4501c1ff9e010bfe26ff5c;
mem[350] = 144'hfb7cfe35025d0110035d0571008dfe7200b5;
mem[351] = 144'hfef0ffb1012a005e037e03d801f500e4fefc;
mem[352] = 144'hffa5ff440083fd7f008bff2aff1dfe7bfdd2;
mem[353] = 144'hfed802c50159fb1ffc64fd9cfdc9003afc55;
mem[354] = 144'h045704440018ff7702a4ff1dffd3ff980483;
mem[355] = 144'h013603ea0097fcdefef10170feb9faa8fae0;
mem[356] = 144'hff2001cb004bfe33ff41ff0dfed4fd13fc43;
mem[357] = 144'h0583066a000700d0fad3022005490523ff82;
mem[358] = 144'h01ee00a8fef200db03ee006dfde6fba9fffe;
mem[359] = 144'h0729fda6fdf6023609310484fe3efaec0545;
mem[360] = 144'hfe9702db0081fd32fe4efe0dffb5fdddfe67;
mem[361] = 144'hfe7d01460009fb2d0008ff14fd6aff3efca5;
mem[362] = 144'h005b00d90145fca0ffc40111fcedfc95fd10;
mem[363] = 144'h0cda0b62035bfd64ff67ffff081309600518;
mem[364] = 144'h01efffbcff790296ff10fe4cfe99fdfafef6;
mem[365] = 144'h00b0fe83fead011efe4f01ab014a014affa5;
mem[366] = 144'hfd9cfefb015afd3afd56fe30fe4cfef5ff31;
mem[367] = 144'hfe37037b025bfead00dbfe6fff680067fd73;
mem[368] = 144'h00eb00c2004cff2b0128ff83feb200b5fdce;
mem[369] = 144'h0080ffe2fed5ff88fe45ff04ff0bfe270000;
mem[370] = 144'hfeb60041fe3cffc5ffff0026febdfe7cffe2;
mem[371] = 144'hfe960031ffbe010a00fefe34fdfbfe92fff9;
mem[372] = 144'h0142fe75fe0e003bffa5ff29fe570101fed9;
mem[373] = 144'hfeb000a3fe94ff6300450142ff10fe26fea2;
mem[374] = 144'hffc5ff70fe77feddfed5fed0fdcefea50078;
mem[375] = 144'hfe90ffda0136ffe0019ffff4feb3ff66008d;
mem[376] = 144'hfe7cff330056fdddfe25fff9000e0130fffa;
mem[377] = 144'hff12002dff9cff58010fffe1ffdeff44ff26;
mem[378] = 144'hffeeffa200b6ff20feadfdd7fdcbfdefffda;
mem[379] = 144'h0063ff46feaa0068ffaaffa300d8009ffe49;
mem[380] = 144'hfe7300df01d40084004c01d60071ff58ffc9;
mem[381] = 144'hffb50087ff6e012e007e011cfee1febdfe4e;
mem[382] = 144'h008afe29ff44fec9ff70fdf0ffd80179fe6d;
mem[383] = 144'hfddbfe3f00fefe4dffc8fedafdd6001e0066;
mem[384] = 144'hfea0fdbbffe0fedd0019ff59fe1fff2efd5f;
mem[385] = 144'hfeb7fd2afe9900620007ff6ffedf0060fd63;
mem[386] = 144'hff05fdabfdc9ff27fdfefe6ffd5900a2fe48;
mem[387] = 144'hff92fe6300c80268ffabffb300d6ff57fed4;
mem[388] = 144'hfe7bffb2ff43023efff1fd98008eff04ffe9;
mem[389] = 144'h00b3ffa8ff24ff7a0087fea60029ff280118;
mem[390] = 144'hfdf9ff3cffdfff8afeadfd3dfd7afd7ffe7b;
mem[391] = 144'hfe6afe80fcc8fe6bfe7afd25fdc600bdfd7d;
mem[392] = 144'hfd8500a4fda8ff5afefbff72ff83ff3ffdc3;
mem[393] = 144'hfda9fe78ff0002f2ff170075fda10094febb;
mem[394] = 144'h005900befdba002cfe92ffd3fd1eff28fe91;
mem[395] = 144'hfea000c3ff73ff83fe96fe12fda2fdc50121;
mem[396] = 144'hfec3feefffcb016501920199010dfec0fefd;
mem[397] = 144'hff19fe3c009d00d8003d01a40152ffd8ffbb;
mem[398] = 144'hff0bffc2004cff37fdd9ff05fd71fd7dfce5;
mem[399] = 144'hfe3cff00fe3a01b3fff200e3fe8f00b5fcd0;
mem[400] = 144'h014b00abffd3fcfaff62fde9026200a6fdb1;
mem[401] = 144'h0014008e0019fdd8ff0afe9c001d014dfbed;
mem[402] = 144'h04ac03c502f5fff10321fea2010e0012015d;
mem[403] = 144'h006a04140293fccb01b4003cff9ffe50fb4f;
mem[404] = 144'h004203a500f2feff008afed200f0ffe3fbbe;
mem[405] = 144'h052203d400150328fecc006d002905faffd6;
mem[406] = 144'h038201650128004d04affeecfff6fb80ff33;
mem[407] = 144'h04aa0138011203c904b004dc0149ff6502f5;
mem[408] = 144'h0161013900e7ffea0054ff4802100026fbf4;
mem[409] = 144'h0380ffc1ffe8fe4500c6ff21fed9ff3afd23;
mem[410] = 144'h01f9021bfff10120006bfe2cff810061fb3e;
mem[411] = 144'h06dc0c590461fd0a01cc0111061b07960355;
mem[412] = 144'h00cbfed900eafe1bfe96fd7c029e02c5ff3c;
mem[413] = 144'h0102009d012f017aff6c01f7fec70119011a;
mem[414] = 144'hffeafe4c015cfeadfe37fea5feed0133ff93;
mem[415] = 144'h027502b4fe9f0090ffd8003600370055fbdf;
mem[416] = 144'hfcf5fdcdffd1fe44ffb1ff3bfc7dff89ff01;
mem[417] = 144'hfd81fcd2fcf8fe57ff80ff8cfe97ffb9ff9a;
mem[418] = 144'hfdc90121fe40fee4fccafe20fee90000febd;
mem[419] = 144'hfe1bfcd2000f00c8fe53ff16fea8fe1600f8;
mem[420] = 144'hfbd8ff69fea8ff89ff68ff8000a5002e004a;
mem[421] = 144'hfc24fd10fcf0ffa0fe45fe47fca3fdcbfedf;
mem[422] = 144'hfd3e00a8000dfbbffe8afe0c00b5fe61ff0e;
mem[423] = 144'hfc85fd62fd54fd1cfdad006e01e4003efd0b;
mem[424] = 144'hfe2bfd27fedcff20ff4dff54fe3efda500a7;
mem[425] = 144'hfdf1fe96fe71fd62ff49fdcbffaffe6d0031;
mem[426] = 144'hfd80ff76ff19fd1efc70ff5dff3c005ffe49;
mem[427] = 144'hfd060062ff4aff1dff1dfdfbfd60fdf6fa94;
mem[428] = 144'hff40fe55014dff230110ff4e0069fe8fff9c;
mem[429] = 144'h01d7012e0054012b018efe3401cdfe600122;
mem[430] = 144'hfef3fe8dffaefdb8ff47fb0afcbcfe72009f;
mem[431] = 144'hfc72000d006ffd8fff16fe50fe5dffc1fd56;
mem[432] = 144'h010300d0fe0000d90149fec100370155ffb5;
mem[433] = 144'hfe8200c4fdce002000c00127ff10feddfeda;
mem[434] = 144'hff65ff5a01cc00040083fec4ff81fe0a0131;
mem[435] = 144'h014000fa008dff75feb9ff3ffed1ff8e003c;
mem[436] = 144'hff57ff9bff2afdf9ff5e0022000efde100db;
mem[437] = 144'h00c6fffafddafef2fe27002b00500045000b;
mem[438] = 144'hfda7005c0069ff6700b9ffceffc100bf010b;
mem[439] = 144'hfdeb0152fee6ff0a01e7003e0218ff12012b;
mem[440] = 144'hff0aff9efe0afdeefe46fde20096ff660115;
mem[441] = 144'h00ef01d40010ffd8fe4100a5007ffe2f004c;
mem[442] = 144'hfedb0092feccfe810170ff58ff17006a00b4;
mem[443] = 144'h0011011d0056fe670018fded004c0146ffbc;
mem[444] = 144'h019f0154ff2aff9e00ff0112ff7e00a10166;
mem[445] = 144'h0149004f0139fe79ff5b01a1fe4700f400be;
mem[446] = 144'hfec7ff220039fea20036005800beffc0fdbf;
mem[447] = 144'h0130fdd3fff5ffe2febcfef5fe46ff50ff7a;
mem[448] = 144'hfee8feb8004e0047ffab0091ff5ffe3efe89;
mem[449] = 144'h00fd0177ffdffea3011ffdd0ff5200dafe94;
mem[450] = 144'hffd4fe82ffa70112ff700165fe480137001e;
mem[451] = 144'hfff4002afe5bff4dfffa00750140fdd8ff3c;
mem[452] = 144'hfe1cfea5fe6a007101320078003efe2effe8;
mem[453] = 144'hfe6700440168ff1a00ea00450071fe1300b5;
mem[454] = 144'h0084fdfdfdf5ff75004100fd008bff62ff50;
mem[455] = 144'hff08fe2000d600b700a9ff50fe73fe72ffb7;
mem[456] = 144'hfecb006afe74feb6fe03fde4fec8014f0059;
mem[457] = 144'hffc80056fe0600930051fe9d005bffd0ff4c;
mem[458] = 144'h00c0ff630025ff30001afdedfffffddcfee8;
mem[459] = 144'h00b30156ff61fdf0007bfe9e0078013fff62;
mem[460] = 144'hff6a0132016e0007ff64fe52feb000befe3b;
mem[461] = 144'h008a011afef6ff5afe2c01e2ffefff740152;
mem[462] = 144'hff8400e4ffd0fe3a0049fe40fe5efee00144;
mem[463] = 144'h011dff2ffef9fe70013dff36ff2aff6600bc;
mem[464] = 144'hff3cff70fb90fa4ffc93fd49fe17032003c8;
mem[465] = 144'hfec5fe67fef6fe26fec8fbc2ff9803b90302;
mem[466] = 144'hfad7fe66fa37f9c2fbd7faa7071605fe01bb;
mem[467] = 144'h000efe5dfcc2fd40feb9fb78ff0902ea02f6;
mem[468] = 144'h00fcfe0e0052fd44fdc8fb25001d02b7fff7;
mem[469] = 144'hfede018b035cfeebf728fc95f957fe7503a9;
mem[470] = 144'hfdc9fdbcfca5fbebfc3dfd3f029200290136;
mem[471] = 144'hf7a8fc49fe74fd25fbb5fd5204bafd07fe74;
mem[472] = 144'hffd0016cffb3fd9cfe02fda3000e030201ff;
mem[473] = 144'h00c000b8fdb9fdd2fb75fd5dfe5e022b02f9;
mem[474] = 144'h014cffad0060fb99fcc9fae2fd5f018b012a;
mem[475] = 144'hf827fee00042fe29fc7ff900084705a6fde7;
mem[476] = 144'hff45fde5fe4c01dafe31ff600071fea9ff4b;
mem[477] = 144'hff9f016d005200c0fe8f0132ff6000bc00dc;
mem[478] = 144'h00bffda0ff7e02e302f2fe4efbb2027b007d;
mem[479] = 144'hfeba01d80018fca0fdbafc11fe9d033801e2;
mem[480] = 144'h00e900f3fa74fb8dfd6dfeee001200630196;
mem[481] = 144'hff7e011efb78fb87fcbffd7500e0ff8bff9a;
mem[482] = 144'hffb8f957f53ff88ef996fe1003ae030d06e3;
mem[483] = 144'h001c008bfbe0ff59fbecfcfc03a4fd72feac;
mem[484] = 144'h015001eafd70ff1afcbcfbf30377fdbc010b;
mem[485] = 144'h07d3044c04adff54fc2bfb2c02e601aa010d;
mem[486] = 144'h0090fd3bfa9cfc68fa1f01a4fb97fc7401e6;
mem[487] = 144'hf9cef7fdfc3dff19fcf10249ff37fc500234;
mem[488] = 144'h01880046fd38fd49fea9fcfe030100d900c5;
mem[489] = 144'h00e70034fe73fcd0fd3bfbbc015dfc250186;
mem[490] = 144'hff2aff06fd8bfa1ffdddfcefff7cff32feec;
mem[491] = 144'h087509d30488fef2fecc00a407ca0b6200cf;
mem[492] = 144'h0184006dfe5f00b10071feacfca0fd680105;
mem[493] = 144'hff43013700d9ff76ff01ff020132010a0067;
mem[494] = 144'h000efedffea5049301dbfedf016b0276fe51;
mem[495] = 144'h0276005dfcfbfdcefd3ffeb801ad00f0fd76;
mem[496] = 144'hfd9ffdccfffb0147ffd7ff02feb1ff69fede;
mem[497] = 144'hffbcfe7bffd40136ffe7fdad014f00eb0152;
mem[498] = 144'h01f20132012200530106ff2afef9fefeff4a;
mem[499] = 144'h00eeffc00088fed500e2ff1eff76fea1010a;
mem[500] = 144'hfe1500860049ff490023ff15010c006dffd3;
mem[501] = 144'hff4b007cfe2bffbf007dfed101f2ff4ffdd7;
mem[502] = 144'h004cfe37fff9ff25003afe3f007efeeb00e0;
mem[503] = 144'h0063fe21fe36ffc8fe0801090178009bfef4;
mem[504] = 144'h0073fdf2ff18ffa7fe7d00f4011dff9300c8;
mem[505] = 144'hfe64012cff290128ffeaff7cfeb6fe9efe42;
mem[506] = 144'hff4cffc7ff460002ff720250fea6fdf4ff7e;
mem[507] = 144'hff22fe23fe35ffaeff1b0056001301cdff47;
mem[508] = 144'h017f00f80142fe76ff42feebfeb60119febd;
mem[509] = 144'h0163ffd100dc01a600fd00b7fe61fe890143;
mem[510] = 144'hfe84ffbcffb70142ffe1ff81ff2400cf0054;
mem[511] = 144'hff88001bff8b002500a3fe720085ff3c0105;
mem[512] = 144'h03e2fc2afb15ff160096ff0e04ccffde0055;
mem[513] = 144'h0318fdeafd60fee4ff26fd1f046602abfdbd;
mem[514] = 144'hfbb3faf2fca0fc41fc03fae203cdfe190266;
mem[515] = 144'h0117fedffd1901b8fe7afaad035a000dfddc;
mem[516] = 144'h02620050fe17ff13fd96fb84025b02caff5b;
mem[517] = 144'h046e01fe01a9ffc0004afb3702de03ae00ca;
mem[518] = 144'h0469ff8efbd9ff77f980fc40fe7ffced0005;
mem[519] = 144'hfc91002b02a4fc72f7effc67ff72fbc1014f;
mem[520] = 144'h01b4fdb6fd29ff9e00bcff170468ff2c0031;
mem[521] = 144'h0373fcf1fb3b0045ff0efb2f05480138fd81;
mem[522] = 144'h0177fdf0fd89fdcdffeffabb008a023bfd9d;
mem[523] = 144'hf4eefd8b0385ff76fcb8ff37051a00c001f5;
mem[524] = 144'hfe68feb5ff28ff83ffca0027fe62ff640098;
mem[525] = 144'h01780032ff5b015ffe50003001d40009fe5a;
mem[526] = 144'h013ffd32fc540485037502b0012c01fffe4a;
mem[527] = 144'h01e5fda0fb92ffd60001ff5d02f30086fd65;
mem[528] = 144'h00e1037403e0011c00a705f702b601b7fdf8;
mem[529] = 144'h01e70308043d0177011b036002a2ffe7fd30;
mem[530] = 144'hfba5fca70cc3ff88f993fe6700ccfe9afabb;
mem[531] = 144'hff7b01fb06c8016000f7012a02e600a0fedf;
mem[532] = 144'h01b002390301014a0028002303d40127fd3a;
mem[533] = 144'hf741fecffd7f04d00539fce7ffcf002bfc8b;
mem[534] = 144'hffc2045605bdfd47fd3a035006c200dd005a;
mem[535] = 144'hfdee02720636ffc0f67ef99c04acfff100a0;
mem[536] = 144'h0054037704d0030c013a02a30341feb10024;
mem[537] = 144'h00d40144016400a60439050b0567fe85fa55;
mem[538] = 144'h02a0002a033000bc01420272051100b5fd13;
mem[539] = 144'hef21f2effcdc021c023602ccf126f512f9d1;
mem[540] = 144'h01ca02db0099fd8c017c0170025c00040018;
mem[541] = 144'h00c1fe24fef0fff100150151fe28ff54fe84;
mem[542] = 144'h04c6035a0450ff6104a7034f002e011703d0;
mem[543] = 144'h01f200c70508004b037703d101ab005cfed8;
mem[544] = 144'hfdaafdd8fefdfee30069fe60011f0097fe6d;
mem[545] = 144'hff99ffe4005efe91009600fd01300048fe34;
mem[546] = 144'hfe25fe76ff2e0084ffb900c2fdb6fe41000c;
mem[547] = 144'h0014fe95fd9efe42fddb0047fe9000bfffd8;
mem[548] = 144'hfe5afee8ff09fda4005bfdeefeacfe900006;
mem[549] = 144'hfee8ff64fe8e003efe38ff63fea7fdc0fe46;
mem[550] = 144'hfee3ff5a009ffdc5ff6cff40004cffa2fdd8;
mem[551] = 144'hfe5f001e0066fec000d6fdcf0064006cff54;
mem[552] = 144'h001dfe15fe8cff13ff5b007afe87feb90094;
mem[553] = 144'hffad00cbfe00ffc1005700e9000afde90013;
mem[554] = 144'hfe2bfea6ff26fe90fef60135ff1200d3fdb9;
mem[555] = 144'hff07fff2ffa00109ff97fe8700a7ff44ff6f;
mem[556] = 144'h002101a6ff3d01170108ff8a0012feac0011;
mem[557] = 144'hfed8ff30ffa3ffffffdfff00013d01bcff22;
mem[558] = 144'hfffbfebdfdeffe4d0066fefefdbf011400eb;
mem[559] = 144'hfe9bfe61ff4e0069ffeffda40120ff8ffdd7;
mem[560] = 144'h05eb05fb006fffa6ff8efe54047404b50387;
mem[561] = 144'h05f9040801870200fe18003c02aa016b021f;
mem[562] = 144'hfe98f869fbad008effa4053cfcb0ff62fb67;
mem[563] = 144'h04c402930364ffb7016e00f50476ff26fd3b;
mem[564] = 144'h064803c6032c00df0020feef02bd004fffa7;
mem[565] = 144'hfae602f2046800c6fee8f765fddcfe7400fa;
mem[566] = 144'h01e002e80293021ffea203c6ffccfebcfcad;
mem[567] = 144'hfa45f7bf01be003effea0534f92cfb9cfb8b;
mem[568] = 144'h03d60470032c01a8002e01a3018b01b800f7;
mem[569] = 144'h06a302ef0317010dfe8bff3f02c6ff520009;
mem[570] = 144'h070c035602d9ff4aff89fff70187002cfed5;
mem[571] = 144'hf569f046fdb400f1fd3a0478f9fafebb0058;
mem[572] = 144'h00c200e5010c0195febfff9dff26fd93ff0d;
mem[573] = 144'h0007fe36fed4ff4aff35ff3f00a3ffccff9d;
mem[574] = 144'h05c60448ffd40090ffccfeef035f0591051f;
mem[575] = 144'h03ca060d024b0150ff4a014f01160291fefe;
mem[576] = 144'h06e9056803b302e5fefeffbc0213050205b3;
mem[577] = 144'h064b03fe028002d0ff720066027505b005f3;
mem[578] = 144'hfc23f8b4f60500cfffddffe3015d04e90331;
mem[579] = 144'h0313033b028affc400690018ff50055000bd;
mem[580] = 144'h05c5068601890149ff3aff3b010104900192;
mem[581] = 144'hfa0f03d90787fc09f69ef5f2fb2501cc033e;
mem[582] = 144'h012d015efdf3ffe4fd110013fbf5fb52fafc;
mem[583] = 144'hf7faf47ffb6efef1ffd1002afa33f763f813;
mem[584] = 144'h06c203f100d0009800b4ff74037906c505b4;
mem[585] = 144'h0369067e029a00930055fea2fd9404d40831;
mem[586] = 144'h03fe04840660ff5afeb4fd09fec001c9023f;
mem[587] = 144'hf74af94001d7007dfd9efd9403860be2ff5a;
mem[588] = 144'hfc9ffef900cc02120047fe41ff2afcc0fd28;
mem[589] = 144'h003b01cb0050ff9800c0008d01a2019e0011;
mem[590] = 144'h02440069005504c2ffae01ea0271069c05de;
mem[591] = 144'h058405cc04c801baffecfdefffc606200519;
mem[592] = 144'hff8fffe601410150ff89fee9fe14fdeffef0;
mem[593] = 144'h0126012700dfff23ff77ff480177fe62001f;
mem[594] = 144'h0007fec700cafee5fe9501260147015f00ec;
mem[595] = 144'hfedc00e4ffa000e4ff14feb6fe030103fecc;
mem[596] = 144'hfe1afeea0026fed6fe48fe7800e800a5005a;
mem[597] = 144'hfe44ff46fddfff59000dff81004ffe57ffec;
mem[598] = 144'h0037fee6fe7100b2ffbdff0e00dc019e00ba;
mem[599] = 144'hfeb3fea8fed40103ffa2fe39ff9ffec10003;
mem[600] = 144'h0031011efdef004dff68004efe1e01530056;
mem[601] = 144'hffb1fdd500fffff3fe64fed5015f0132ff43;
mem[602] = 144'h0018fe1afdf3022c00000034fef2fe17ffae;
mem[603] = 144'h010100490061014b0000fe23fecc0125ff43;
mem[604] = 144'hfeffff85ffd500210147ff09ff5b0050fe7a;
mem[605] = 144'h00c7009bfec100daffd7fe37fea7fe7201d5;
mem[606] = 144'hffd4fdb5feecfed5feb40161ff2fffd200e1;
mem[607] = 144'h010e007c0005007bfdbefdb5feb3fde500f0;
mem[608] = 144'hfee800750039fb67febd0165ffd8fd0dfc6c;
mem[609] = 144'hff5a0103ff1efc5c003c016eff32fd11fc67;
mem[610] = 144'h02c507710a27fdc70015009efefbfb71f9a9;
mem[611] = 144'hfe4001cf034ffbacff23fe90ff12fdc2ff9c;
mem[612] = 144'hfdb701320001fe93fcf200ddff2dfde3fe93;
mem[613] = 144'hfc18fd43fe0d0352fbb300d901eafdb6fc5e;
mem[614] = 144'h015f03ea04bcfd64ffcbffd9028705a50463;
mem[615] = 144'h094d0bce0a1ffcb4029903bf05d20317050e;
mem[616] = 144'hff44fe270279fbd3fe0b0074fddaffc1fd4e;
mem[617] = 144'hff38ffa5ff91fc2dfe1dfffa002afee4fdb0;
mem[618] = 144'hfd6c007afffbfc70ffb200a4ff56ffabfdca;
mem[619] = 144'hf8cdf553fbbe002c01c40123f4e4f76cfa9a;
mem[620] = 144'hfea101bcffd7fe7aff67005b0166fe7900cb;
mem[621] = 144'hfef7fe740157ffabff08fef10078fe2d00a1;
mem[622] = 144'h027203da0007ff9ffe56028600a7fe850065;
mem[623] = 144'hfe0200bdfee0fba40045013bff77fff0fe5c;
mem[624] = 144'hffcaffc6fe13fe060199fff40151ff33016f;
mem[625] = 144'hfe4a012fff3a00d10001fdd6ffaffe250080;
mem[626] = 144'h00bbff8affb0feb9fed80131020dfe9effe0;
mem[627] = 144'hff4a0198feaa012efe750077ff5ffdc8ff20;
mem[628] = 144'hfeceff1afef3000aff54fe4fffa0ff16fe1b;
mem[629] = 144'h0027001bffb5fe9fff0cff0700a9012f0100;
mem[630] = 144'h01f200f4011d0185001e0114fdbfff6300d9;
mem[631] = 144'hff9cff00fe5eff2d001bfecb00010067ff39;
mem[632] = 144'hffa70119014a00cf00a5fec2008cff05ffdc;
mem[633] = 144'h01aeff7200380123014f00effe8afe81ff2e;
mem[634] = 144'h003b0044005f009e011bfe76fff7ff220002;
mem[635] = 144'hfea500a3ffabffbaff1dfe87fdd4ff18ff88;
mem[636] = 144'hfff5fe5600b6006dfeb7ffec014f01260145;
mem[637] = 144'h017b00bbff8c0063ff3bff7301b1fe24fe4c;
mem[638] = 144'hfeeffe34fefcff23fe0f00190112ff320119;
mem[639] = 144'hfde201760128fde4fe86ff7d00ce015dfe36;
mem[640] = 144'h034a02060293f847f960f993020bffcefdb0;
mem[641] = 144'h0304011c00c0f907fae7f93affbe0156fedb;
mem[642] = 144'h005dfd1af91ef759fe01040702e0feec0462;
mem[643] = 144'h01ab025a0289fab7fb95fc57ff8dfe4efcba;
mem[644] = 144'h032401700291fcf1fcf0fd4400a1fe56fc0a;
mem[645] = 144'h055a0327033c0033f5a3f46a047a012cffac;
mem[646] = 144'h030afd21fdf6fb5a02920228fcccfc24ff6f;
mem[647] = 144'hfdadfa92fc28fe4e07140c48fc97ff8affe7;
mem[648] = 144'h019d03390251f839f9d4fba200d8fe68fd2e;
mem[649] = 144'h04d70149027ffadcfb0ef8dd019cff05fde1;
mem[650] = 144'h029d04b90273f9e7f9abfab4ffbdfe68fa98;
mem[651] = 144'h036a0bec0568f93cf9eb011c02d004a201b0;
mem[652] = 144'hff4f0011ffdf01cffe3ffeb4feecfe5c0067;
mem[653] = 144'hff6fff950000feea0010017600f2fe20ff8c;
mem[654] = 144'h01db0138ffbd026ffd9afb3201ea00ca02dc;
mem[655] = 144'h04d802a7024afb28f8b7fa74020b00fcfbe0;
mem[656] = 144'hffdcff2efedb0029ff4dff62010900560007;
mem[657] = 144'h0073fe98fe0d00680180013bff0dffce0064;
mem[658] = 144'h0017ff5eff240146014001b3ff97ff9c0149;
mem[659] = 144'hffe3ff5700fbff4f002700d30138014b007f;
mem[660] = 144'hfddcfef601520028fe2bffb7014dffa3fea3;
mem[661] = 144'hff32fe90fe11fe44ffedff07fe5dfe0ffed2;
mem[662] = 144'h0054ff88ffcc0024011d0161ff8dff5a00fa;
mem[663] = 144'hff6e012cff31ffa5fe0ffda5ff4901f30193;
mem[664] = 144'h00b7fff9005c0009feca014cfe18001f007b;
mem[665] = 144'h0141fee9ff72fe40000dfeadffd1fe4200bd;
mem[666] = 144'hffb4ff9afda80097feeafe4c01b200b10061;
mem[667] = 144'h001ffeb5009001dc011d0006fdb000250097;
mem[668] = 144'h00caff58ff46fe440182ff0ffe2800d1ff65;
mem[669] = 144'hff73fed90006fe7b01ceff5100aeff95fef4;
mem[670] = 144'h0079ff55ff42ff400118ff36fef2ff80fffc;
mem[671] = 144'hff620095ff95015d00bf003efdc8fe7afffd;
mem[672] = 144'h043f0130ff6aff20ff05fea800c90221fefc;
mem[673] = 144'h053203e7fe9cff6f0116002d0272042bfe9b;
mem[674] = 144'h019100fcfe04fd92033601730224fda80123;
mem[675] = 144'h044e0441ff2dfd57fec4fda3ff2c00ebfc98;
mem[676] = 144'h05f004bbff7400ad00b1fd71007d0175fd2c;
mem[677] = 144'h011505e401f3ff6bf705fe0efcf803100138;
mem[678] = 144'h061cffd4fb9200cb0357fc89fddffc6d00c7;
mem[679] = 144'h0480ff25fd8dff7d07d6026bfc90fd9f0285;
mem[680] = 144'h04b1016400f8fe7a00ebfe6f0312015ffe65;
mem[681] = 144'h0455031f010d000bfcdffb34fec30392fb05;
mem[682] = 144'h05ef04ba00440233003eff52febf02b0fd61;
mem[683] = 144'h034b003c02f1fbacffcefeed0684fadc006d;
mem[684] = 144'hffd3fe7201a0007200c5016202eb01d3ff3d;
mem[685] = 144'h0074fee2017101a700e10012fecb00c700e9;
mem[686] = 144'h02d4030300490266ff7a00a9053c02a0005c;
mem[687] = 144'h04dc03fa00deff69ffe2fd6a0203043efbfb;
mem[688] = 144'h03540007f90cff49fd0fff0701c8011b008a;
mem[689] = 144'h01290016fbdffe4bfe51fbed00f800da01c5;
mem[690] = 144'hfcdaf592eed7fe96fcec007d067102d2fc3d;
mem[691] = 144'h0380fcf4fb1b0128006dfdc002e20228010a;
mem[692] = 144'h0282fee4fe73fef4fd7afb8102ca047b0250;
mem[693] = 144'h07d501c50286002305ecf6f0002c004c030d;
mem[694] = 144'hff1dfca8fc6fff25fcf902f10317014effcf;
mem[695] = 144'hf5acfe09fec4ff360076046e0695ffa8fe85;
mem[696] = 144'h00a8ffb8fab6fdfdffdcff0c034603450083;
mem[697] = 144'h0338fe89fa00fff8ffcbf9de0401034502c1;
mem[698] = 144'h02bb00acfc67ffd9fcd0fd1a041203d6012f;
mem[699] = 144'hf9b0fb8d00d00016fe9fff01029e07d60556;
mem[700] = 144'h0019fd56fdb30183011dfe6cfe41fd960117;
mem[701] = 144'h001e018cfe8c0131010d00d8001901270194;
mem[702] = 144'h029dfe68fc700055009ffad9005c01c3fef3;
mem[703] = 144'h02cf002ffb4bfd41fc49fef3030700e4ffdc;
mem[704] = 144'hfddcfe55fba0016f028901c0feea011f005b;
mem[705] = 144'hff27fddcfcc8fdab0257026efdbd01ca00f8;
mem[706] = 144'hfb010061fd810235041b006a052503a5fbdb;
mem[707] = 144'hfe77fcaffed2ff4a00e7fff8028702e7ff8d;
mem[708] = 144'hfdd9ffd7ffd2fdbd0285014c005b03460087;
mem[709] = 144'hfe5bfeb8fe01fcb30151fec8f986ff1e01fb;
mem[710] = 144'hfd18ffb600be024002550375082c015cff01;
mem[711] = 144'hf89bff12ff2b0248ff1d003809f2017efe50;
mem[712] = 144'h004ffd0bfcb100dc0269019e00f80064ff09;
mem[713] = 144'hffb8fe45fee7fd9a02b90194fe85036fff5c;
mem[714] = 144'hfdf6fd3ffdabffa0037f049a03ee04110185;
mem[715] = 144'hfdde00c8fc7d03fd0291f7a4ff7c0050ff78;
mem[716] = 144'hfdb8002f010f00d1024ffe69ff8e006e00a9;
mem[717] = 144'hfe96fec8011dff5afe29011d019901c5ff68;
mem[718] = 144'h0244fd13fee2ffcf011efdfcfb98fec9ff7a;
mem[719] = 144'hff90ffc5fd66fe4702c700770021010bfea8;
mem[720] = 144'hfef002140773fe9eff1d02a7007ffd5afe78;
mem[721] = 144'h01dd01ff047100d30091ff3401beff11fff6;
mem[722] = 144'h0084fdec09f0fe7ef7d3ff2efe4300830017;
mem[723] = 144'hff7c01b5067e02b9ff8bfd96ff42fd63fffa;
mem[724] = 144'h000401d40477ffd6fe4bfed80104007cfdd7;
mem[725] = 144'hff00fe4efec702f8fe920085058afeedfce4;
mem[726] = 144'h022f03390364fc6ff910ffd1fff2008c0158;
mem[727] = 144'h0198015003e8fd85f900fc7bfdec0291021a;
mem[728] = 144'h025c00ec064e011ffe9f01590258fdb1006c;
mem[729] = 144'hff72016403b601c500a8004c0427fce5fd4c;
mem[730] = 144'h028f015103eaff14fe84ff62018efdebfd06;
mem[731] = 144'hf765fd96fe880077ffc40200f7be0226fc6b;
mem[732] = 144'h004fff2b0264ff5a0039002b02b8ffef026a;
mem[733] = 144'h01b8003600f200fc007bffe0feb4fea2ffce;
mem[734] = 144'h029903ff04b0016e06b503bb03a6feba044b;
mem[735] = 144'h023302d1036901ceffdeffc102a6ff38ffb7;
mem[736] = 144'hfe2efe7efe110182ffdeffb4003200cdff97;
mem[737] = 144'hfdbe00e10142010bfe6aff48013dfe5ffdbc;
mem[738] = 144'h018801d7fef4000f007d003aff26ffaf0109;
mem[739] = 144'h0140011100c5007dfe810098fdbefdecfea7;
mem[740] = 144'hfe4dfe970075009a00d3ff940078ffc3fedf;
mem[741] = 144'hffd800bbffcd005901730098ff87fdce00f7;
mem[742] = 144'h010dfff20059fddd00d4fe5700f1feb1ff08;
mem[743] = 144'hfe5a016a014600e2fec4fdcafe58018c002a;
mem[744] = 144'h00f1fefbfe4200b5feb000f5fdcaffad0105;
mem[745] = 144'h00da001600fc01a5fe6900e3ff790058ff3f;
mem[746] = 144'h00a6feacff3a0034ffb2ff41fe18ff81fe88;
mem[747] = 144'hff38fe8b0011ff4800cdffbefe77ffa1000a;
mem[748] = 144'hfef0009701b800ba005f0147fedbfe24fe2e;
mem[749] = 144'hfe4a0139ff0200f6ffd1017e000cfe27feb8;
mem[750] = 144'h00bafec9ff840083ffd3ff2f0065ff1affb3;
mem[751] = 144'hfe10ff9301150126ff5a0131ff7b017cffa5;
mem[752] = 144'hffccfe6101bbfaa2fab6fc63ffe7fd2afd4c;
mem[753] = 144'hff31ffd9012efb9ffad3fdbe01830017fbc6;
mem[754] = 144'h00a5047c09c5f648fab5026d010e00c901fe;
mem[755] = 144'h00c801220264fabafc86fb4d026aff22fc3d;
mem[756] = 144'hfe17ffed024afa57fb21fc1800cafddefec5;
mem[757] = 144'h0394fef1fe760028f5edf98d049dfe4dfe50;
mem[758] = 144'hffb3ffcb0125fb9ffedc01ec0167fe9700e7;
mem[759] = 144'h054c01410120fc23fce009d001fb05ca063e;
mem[760] = 144'hff67015b0089f8d2faddff080133feaefbd3;
mem[761] = 144'hff3101e7016efa79f98dfe9a01c5ffccfb70;
mem[762] = 144'hfe2d004700d7f7b3fa07fe1101adfdabfb6e;
mem[763] = 144'h05d50a0d0118fb8efabcfe1dff62fe10fd3d;
mem[764] = 144'h003f00d1fef00180fec9fee202db002d0011;
mem[765] = 144'hffd4001f0134ff38fff3012fff3e009dff76;
mem[766] = 144'h00ab00d2042402effdcafe2e0231015bff5b;
mem[767] = 144'hff0bfef70198f8e9fba4fe4500cffd7dfdd4;
mem[768] = 144'h000fff88fd4ffd0dfeeef8ccfdcb027702df;
mem[769] = 144'hff55018cfe20fe54fd91fc94fdca0356ff9f;
mem[770] = 144'h01f30309f599fe3affc9fc990617030808f6;
mem[771] = 144'h02ac023fff42fff6fde9fc2dfb18ff61ffac;
mem[772] = 144'h00a700b8fd36ffb400dcfa58fdc2000301a9;
mem[773] = 144'h041e031003befd17f7c0025e000004a7017a;
mem[774] = 144'h01e20084fbceff5d0208fb23fa6dfc890297;
mem[775] = 144'h01a400a6fc8200d2048c04280057fbbb059e;
mem[776] = 144'h02a4ff38fd1afe1ffff0fbd5006c025800f5;
mem[777] = 144'h021f0199fe09febdfdc2f93bfd5a003d02b5;
mem[778] = 144'h019a01eeff4aff09fde2fb3ffb8ffe9d00f8;
mem[779] = 144'h06fc0d2004dbfdf3fe36fa5b0e150da00645;
mem[780] = 144'hffebff64fef7ffc7007a0066ffdcfe3dfe51;
mem[781] = 144'hfe21fe42fea1019c01c8feaeffa20161fe74;
mem[782] = 144'h0069fddfffb000d8005a01070000011bfefc;
mem[783] = 144'h0210ff9400a5ff58fe9ffadafdaf01e502a2;
mem[784] = 144'hfec7fe64fdb0fe85ffb1028e0083fd7ffe9d;
mem[785] = 144'hffc0fe37ff74feec006002ad040d0086ff23;
mem[786] = 144'hfe6cfeb7036dff7cff1c03b30530ff82fbd8;
mem[787] = 144'hfd9dfed4fe5ffd5dfd2a012e06220248015b;
mem[788] = 144'hfd58ffb000e8fe76fe9e0381051900afffcd;
mem[789] = 144'h051200dcfe35011f0512f907021dffa7ffab;
mem[790] = 144'hfc6400ec0426fe47fe7e08d905be042900a5;
mem[791] = 144'hfd2e030a02b200b1ff9b0499093a05bf0095;
mem[792] = 144'hffe5002fffc3ff68ffd5023102f40128ff33;
mem[793] = 144'h006cfc92fec3fdd50054022e05630000fdd1;
mem[794] = 144'hfcf7fe0afcfbfca5fe2c00600457013afd7a;
mem[795] = 144'hfdc6ff52ff640121ff970329f6d9f891fc1b;
mem[796] = 144'hfdc1fe3e0197ff5d0066fe3fff280100025c;
mem[797] = 144'h016e0011ff6e01aa0159ff8dff14fe5d001b;
mem[798] = 144'h023efe73ff80fe4afedcfcbd0090ff040096;
mem[799] = 144'h011dff93fdc8fe08fef7012a022e0049fcbf;
mem[800] = 144'hfeacfdd4000dff3f009701a5fd9effe90142;
mem[801] = 144'h00daff4fff9dff250024003e00f1fe32fdbd;
mem[802] = 144'hff4dfe0b0117fe9d008800b6ff30ff70fe9d;
mem[803] = 144'hfdef0033fe1cff28ff5dfde1ffc100b4fe10;
mem[804] = 144'hfe6dfe6dffac00effef2ff0fff13fe5f002b;
mem[805] = 144'hfddc00e50020ffcf00effe15ff75fd630076;
mem[806] = 144'hfe4bfe1bfd9eff5ffea1fef80138ff6bfecc;
mem[807] = 144'h01220144fee20075ff12ff38006afe820085;
mem[808] = 144'hff85fdd7014ffe22010bfd3efde200affefa;
mem[809] = 144'h00c6ff73007a00970065ffcffd56ff77005b;
mem[810] = 144'hfdd2fec3fd960124ffeefe2601aefe9dfead;
mem[811] = 144'hffb4fe4efde30091003b00abfd580010ff47;
mem[812] = 144'hffa4ff5000b00193febcffcb000f007001b3;
mem[813] = 144'hfec900fe00ee008fff10fe28fe9b0092ff8c;
mem[814] = 144'hffc40090fffafec0004f006bff09fff8fe1d;
mem[815] = 144'hfd720088ffb7fdd300cffe18ff96fec5fff5;
mem[816] = 144'h0106fd84fb530075fd57fc8a0576046000a2;
mem[817] = 144'h0171fd2dfd4700e1fd8dfba6048c01de012c;
mem[818] = 144'h05c603dcfef3fc65ffa403c20330feb701be;
mem[819] = 144'h037cff0bfd1201affec8fd2b00c9025f047f;
mem[820] = 144'h04d1fe60ffcd0136fd1eff0a014002d500eb;
mem[821] = 144'h09ed005a0065003103aaf79dff4e00890317;
mem[822] = 144'h02f7ff4f0205fe9200d7fe97ff2f051603d1;
mem[823] = 144'h05e0090502c8ff8e00b10613fd1e06f8059c;
mem[824] = 144'h0221ffd7fe0d00e8fe6afe3b03ea022f01fb;
mem[825] = 144'h0403fdf8fc6703d4feddfb9f039004050000;
mem[826] = 144'h02770050fcdf0034fe81fadafff4010e0302;
mem[827] = 144'hfe4d010d01f1fe8afc67090d01fdf57c0001;
mem[828] = 144'hff35feebfebaff32fe1f009e0274fff5ff51;
mem[829] = 144'hff9efe70fe7e004701800000fe4e000dfe24;
mem[830] = 144'hffe1fdacfee60487fe9e00a6043f0098feaa;
mem[831] = 144'h029dfe5afc42022cfc2cfefe038201d10110;
mem[832] = 144'hfeca0256fe68089e03f70467018d020006e0;
mem[833] = 144'h01f8ffd8fee9058806bf0388008801220664;
mem[834] = 144'h0077f8d1f8ff0a2efe4dfc42ff3506180024;
mem[835] = 144'h001dfff7ffdd076906770297020102850678;
mem[836] = 144'h0143009100db0581062203b80324036307ae;
mem[837] = 144'hfe24ff410004ff940ec905c70190fe5a041d;
mem[838] = 144'h00a2031ffed10420fd34fbf3ffe9068d014c;
mem[839] = 144'hfbc7ff3000be03d8f55ef523fd58fef6fb56;
mem[840] = 144'h006c0246ff24078d0650039702b9046a0720;
mem[841] = 144'hfe98fe3d00590648047c053c04cb016008d1;
mem[842] = 144'h015900effea207a20611038603dd03cc055d;
mem[843] = 144'hf9dff8affe2a04ca03b80361ff6e0502fed6;
mem[844] = 144'h0167007900e1ff32fca1ff57ffd2fc3cff6a;
mem[845] = 144'hfeaafffffe8f00fafe5a017901780023feb8;
mem[846] = 144'hff04fe67ff15ff23055c037f011800f90151;
mem[847] = 144'h021e020200f106ae03a202f10045038f0562;
mem[848] = 144'hfcc4ff87024900140055fefdfd09fda8fd8b;
mem[849] = 144'hfe06fe9f04a7035700860078fc5afc4bff89;
mem[850] = 144'h05cb06800fdeff0e019dfec3fab4fb0d0235;
mem[851] = 144'h016f01ea0210032a0064001df937fe32ffe2;
mem[852] = 144'h00f0ff3f041101370229ff50fb09fbf901a6;
mem[853] = 144'hfb52fcb6fc0300c0fb0d0857fee8fd98fb8f;
mem[854] = 144'h05ea016d0565fe6f0017fc81fb280374051a;
mem[855] = 144'h0cd10c8a06b8018b016ffe41faff05bb0457;
mem[856] = 144'hff03fdd7054d013a00a8fe2bfec3fe8e01d4;
mem[857] = 144'hfc41ff25035a0216fff1ff03fe25ffc0fe60;
mem[858] = 144'h0274fef802ca005a01f4ff9ffb7dfce301bc;
mem[859] = 144'hfd2af4b3fd01010b0337ff54fe18eec8fec3;
mem[860] = 144'h00b8ffcf011aff12fff3018a0162019aff31;
mem[861] = 144'h014e01c6013e0060ffb7fee80119fe6ffe77;
mem[862] = 144'hff01006c022f02d4013204660203ff1e0100;
mem[863] = 144'hfe14ff93041e00a00277fec6fd73fe5200c2;
mem[864] = 144'h02da007301a3fe6bfe25ffecfc7300a80148;
mem[865] = 144'h02c002420260fd72ff8a0148fcadfdf3025d;
mem[866] = 144'h005b00c50275fe84059efe3ffbe5fb7d0797;
mem[867] = 144'h005b02ed028afefe00ad01ddfa1cfc0cfe50;
mem[868] = 144'h0292025700adfce2fff7015bfab1fd0a01d9;
mem[869] = 144'h002e026a0291ffc7f8720606031800bcff0c;
mem[870] = 144'h015105460203027c05f1fefef684fa20ff52;
mem[871] = 144'h002804040046014d0a830024faf6fa260162;
mem[872] = 144'h031b02670043ff8a01b7fdcafca3fefe0366;
mem[873] = 144'h02ea03ca03e5fb66fdb6feeafb82fd340256;
mem[874] = 144'h0384000f02e0ff150151ff33f841faea010b;
mem[875] = 144'h011601bb0040fdb900e9fb6805ed05bb096d;
mem[876] = 144'hfff102cafee2fec600d8fe95ffee0048ffd9;
mem[877] = 144'h00880075003e004ffebfff1100baffacfeb3;
mem[878] = 144'h012c019c0219ff79fc2a01b6fe4200bf00c0;
mem[879] = 144'h015700e902aafeec0198ff29fab2fcb302fb;
mem[880] = 144'h01e4035c01f0fac9f9edfaa6fc5f01480008;
mem[881] = 144'hfefb015a01fcfce2f8f6f98dfc9fffb00090;
mem[882] = 144'hfb18fd2df8fcfa99025fff25021901c3ff95;
mem[883] = 144'hfe3500a6fe84fb0afceffb0afbc7fd63fa18;
mem[884] = 144'h005802550015fe07fd5dfe8dfbc8ff5dfed0;
mem[885] = 144'hfca3029c013f003df6dffde0fcd2fedeffd1;
mem[886] = 144'hfe64fdfeff98fd7102ff006dfd65fd99fc75;
mem[887] = 144'hf8b5fa2dfe2ffe6206f7057f01b6fccdfedc;
mem[888] = 144'hffae0315fe02fb3ffcf5fc55fae1005b001c;
mem[889] = 144'h002401b0ff69fa11fbe9fb79f8d0016d0037;
mem[890] = 144'hffb9ff620264fcd1fd47feb2f99effadfe7e;
mem[891] = 144'h02630401006ffb96fe72f79a062d08470274;
mem[892] = 144'h0042feedff2801c001040008fecfff8201b1;
mem[893] = 144'hfe6a01610182fed101d901dbfee2ffb600d7;
mem[894] = 144'h02a5001d00dffd48fe01fb68fe4d01d8011f;
mem[895] = 144'h013e02b20143fd03fb49fb63fde8ff0bfe9a;
mem[896] = 144'h0188034603cc007b00d8026f0018fda4018c;
mem[897] = 144'h01e40077040e021300460073000dff8800f3;
mem[898] = 144'h0020ff710c0effb8fbc9fef0fe05fbccf77f;
mem[899] = 144'h04ed03c606e90237030300b7fdb6ff14fe73;
mem[900] = 144'h0457016703ca0321ffa9fe0cff9ffdf6fdf6;
mem[901] = 144'hfaf1fd8dff9e04b00778fe6b0513fde6fc02;
mem[902] = 144'h030a042b08ae00ceff38f983ffbe00a90077;
mem[903] = 144'h07960944096afee3facff9ebfab4ff02fef6;
mem[904] = 144'h034d039e06a701dd01be003c0227008f01d0;
mem[905] = 144'h02f4ff9a04dd03d70006018801d3fe6efff2;
mem[906] = 144'h0449026a035002d100fdfbab002f00fbfc9c;
mem[907] = 144'hf0a2ef7afadd00f9018305cff7dff7ee0003;
mem[908] = 144'h005e022aff050056fee1002e009f00a1ffd5;
mem[909] = 144'hff6c010ffe77ff0a013afefefe35fe66ff2e;
mem[910] = 144'h016c03db0433006f004c04b10255fefc021a;
mem[911] = 144'h02c2021d053a011e0187ffd4ff580012fde2;
mem[912] = 144'hfd9bfdd2fe84fdaf00f3ffaefd9500fefdc5;
mem[913] = 144'hffb0fda7003cfdfd0000ff5afdb1ff770053;
mem[914] = 144'hfea9fe0c00190078000000baff01ffdefdcb;
mem[915] = 144'hff58ff800080fd7ffe160030fe65fdaffe38;
mem[916] = 144'hff9cfde8ff79fdf900b6ff6efdd7ff68004e;
mem[917] = 144'hfff8fde2fe76fea8ffa4010cfe8c00f7feac;
mem[918] = 144'h006afec9fe4afee0fdc300fcfe37fda70033;
mem[919] = 144'h009cfe13ff88fe2eff78011c01a3ff49ff5d;
mem[920] = 144'hfe5bfe4fff9cffb7fdc40017fda2000f0072;
mem[921] = 144'hfe73fdc20116fdebfff4ff5e009dfd9fffa4;
mem[922] = 144'hfed1fedfff87fe4100c5fdfd0095fded00d0;
mem[923] = 144'hfe52fd8e00b1fdd7fe0efde8ff5c006ffe51;
mem[924] = 144'h0048ff8b0096feadfe6100da003fffbdff8a;
mem[925] = 144'h0157ffaffefa01c700de0160000effd0011d;
mem[926] = 144'hfdc8ff5400170109fe0cfdc800d100fbff2a;
mem[927] = 144'h0063fe0ffe6fffc2fea0fec50043ffdcffd8;
mem[928] = 144'h013202ce00a202e0037a04a2001e0286064d;
mem[929] = 144'h019302bf0179022104b80281006102d0048e;
mem[930] = 144'hfa7dff2afd1e05010013f87102010bd00005;
mem[931] = 144'h00cb003f031005bc05b0fe7100eb061f0386;
mem[932] = 144'hfec402570365019c044c00f200a6052e02c4;
mem[933] = 144'hf6d3022d00d7fea100c606c5f96301db02a7;
mem[934] = 144'hfff70290ff0c0065facffd15053afe2700c9;
mem[935] = 144'hf822f8b9fdf9011cf82af4920239fb3bfa86;
mem[936] = 144'hfe9503a4028104a7059fffb8027d061705ea;
mem[937] = 144'hfeee0401022b01a004c90479ffa8028f0288;
mem[938] = 144'hfefa03b8030402ea02a60078fe3a03a105e9;
mem[939] = 144'hfccf0355017c02850192fb74016b0994fe2e;
mem[940] = 144'hfdaf0107fe5aff1ffcf0ffb0febafee2fed6;
mem[941] = 144'hff8dfe3b017a00f2ff27fea6fe9400edffbe;
mem[942] = 144'hfecf00f6023c02f5050b0553fcb9025c05fe;
mem[943] = 144'hfe6b0162038c02d306f802be00d4040704cc;
mem[944] = 144'h0075ff5e00cdff46fdc60086fda4fd80fd83;
mem[945] = 144'hfef7fdeffd94fe86ff0b00e9ff73fe6f009f;
mem[946] = 144'h0067fe05fecffe25fdfe013800eafe4bffcd;
mem[947] = 144'h0034fda100d800920046fdaf0043ffeffe7a;
mem[948] = 144'hfe52ffd40031fe73ff56ffd6ffc5ffe7000a;
mem[949] = 144'hfffdfea3ff2400c1ffe70021fe0a009000a6;
mem[950] = 144'hfecfff23fd8f007d00ebfd71feaffed6fe40;
mem[951] = 144'hff12ffc4001bfe5bfe37fd9d00cafddcfdd0;
mem[952] = 144'h00f1fe54fd8dfd6ffff00098ffeeff87fdf6;
mem[953] = 144'hfeb4fe1700310019fed0fdbbffaffe94fea3;
mem[954] = 144'hfdbc008dfe05fe0dffaffed9fdf20041000f;
mem[955] = 144'hfe4dfff9ff3800ef002f0094ff13fdb7fdc8;
mem[956] = 144'h014b0173fe91feb4feb500710151004d0016;
mem[957] = 144'hff96ff270066fe27ffef00c6013d0021fe67;
mem[958] = 144'hfe7ffe76fe0efe6ffd610054ff36fed9ff27;
mem[959] = 144'hffce00e0fd87ffadfdefff7efe4efdcfff33;
mem[960] = 144'h00800044fe58fec40112feb0ff97ff31fe1c;
mem[961] = 144'hfef9011fffe700acff6bffc8003301420141;
mem[962] = 144'hfefc01c8005afe39fe010152ff1afe04005a;
mem[963] = 144'h00dd002000f40063fee300a2fee3ffaffdec;
mem[964] = 144'hffebfe9f000afe4cffacffbffe51ff3efeb9;
mem[965] = 144'hffdb0105013bfecb0064fecffff00124ff85;
mem[966] = 144'h013eff2d0133fe63fdc7fe17000d00520069;
mem[967] = 144'h0080ff98ff77003200b100dffe62ff6400d6;
mem[968] = 144'hff5fff9c0143008f00d7ffb6fe6dfe9dff3d;
mem[969] = 144'h00cfffdbfef6ff580088fe3aff59014d0153;
mem[970] = 144'h015d01240118fddaff080180ff02fdddfebb;
mem[971] = 144'hffc3feebff240023fdf900c1006401bf000d;
mem[972] = 144'h00b2ff64ff5100edfeb9fe8c0191feabffc6;
mem[973] = 144'h00ca00d2006c0005fe9bfeac00b5ff5effe4;
mem[974] = 144'hfe3cfe3effe4ff03011800960110fe59ff89;
mem[975] = 144'hfee80009fe66ffc4ff9afdc700d000a8ff48;
mem[976] = 144'hfe0dfe4efec70219fd41fe34feeafda8ff1e;
mem[977] = 144'hfd8afe74fe97ffd2fe30ff5bfdcdfed4fe9e;
mem[978] = 144'hffba02de01d200b0fcb6ff7cffce005400b6;
mem[979] = 144'hfe5bfcc9fe6dffe1ff32fd33006d01f4ff00;
mem[980] = 144'hfe5efd29fcdeffc8fdd7fefdfd72ffb8fe58;
mem[981] = 144'hffabfff6ff7dfcf6027a01e2fe47fec70092;
mem[982] = 144'h006ffe51fce1fcd0ff35fd2aff9200c3fd9d;
mem[983] = 144'hfcbc02f7ff4affeafe5aff4a01d0ffadfd1d;
mem[984] = 144'hfdd0fd92fe0d00e2fe260062ff8bfedf0024;
mem[985] = 144'hfd39fcc5fca0009dffe9fe5afe89fd98002f;
mem[986] = 144'hfd90fcbafd2b00ecffbdfd1afd19fd80014c;
mem[987] = 144'h00100204fdd3ffeafdd5ff9d0013fe7ffd7c;
mem[988] = 144'h008601b700ab01c101aa01480073016e0004;
mem[989] = 144'h01d101d2011401acfeb40099ffe701040178;
mem[990] = 144'h0015fef5fcda0000fd1e0071fe12fd21fccb;
mem[991] = 144'hfe7aff270006004ffc93ff66fd9dfd9cff64;
mem[992] = 144'hfe64fe77fb00fbb9fe2ffe9400cb004bfc10;
mem[993] = 144'hfdc2fd6cfc67fd6cfb14ff5c000bfe88fdad;
mem[994] = 144'h018e0370fcaffee402340408057afd6b0181;
mem[995] = 144'hfc0afd6efd3ffd25fb82ff3402db002ffd6f;
mem[996] = 144'hffa8fefffbedfe66ff6afeb7048bffb9ff84;
mem[997] = 144'h0f0a049501970050fec1fcb1048504d9fe08;
mem[998] = 144'hff33fe4dfdb0014e035906a2013cfe620024;
mem[999] = 144'h009d0088ff0bfffb06ba07d205ed02330375;
mem[1000] = 144'hfed5fe94fc41feaffe00ff260013008afdc0;
mem[1001] = 144'hfdd3fee0f9d6ffa7febaff99ff6f0165fd4c;
mem[1002] = 144'hfccffe29faccfc23fe7502580434ff04fee3;
mem[1003] = 144'h124e11ab04b8fba600ca006606a100aa0334;
mem[1004] = 144'hfff6fec0ffbd016201d5fe5700bc01b90055;
mem[1005] = 144'hfeeaff19018100c4ff87fea800bbfe4200fa;
mem[1006] = 144'hfc19fc8bfcdafe9dfd46fabaff48ff55fc4d;
mem[1007] = 144'hff21feeefd33fc4ffe2bffb902fcff10fc6a;
mem[1008] = 144'h028afee600e401e30274fddafdcbfee2faae;
mem[1009] = 144'h029f00fbff9500340239012effafff29faee;
mem[1010] = 144'hfb67fa3800ae008400e5fcb102f5fef0f7ea;
mem[1011] = 144'h030d008efd5f010300d3fdaffcef00cafd7b;
mem[1012] = 144'h00eaff89feea025602c6ff6cffe1001bfef8;
mem[1013] = 144'hf729ff92ff030350055103dafe860084ff0e;
mem[1014] = 144'h027fff37ff060262feb4fc010160067800fa;
mem[1015] = 144'hff6a006d00dafff6000efc3c02f0010a01b9;
mem[1016] = 144'h01680186ff32ff84ffd2feb4fdd4fe9afce7;
mem[1017] = 144'h01d40133fd8400cbfeabffa1010a02cafb26;
mem[1018] = 144'h0259ff06fdd7ffa70133fddffd4d00ebfdfd;
mem[1019] = 144'hece7e9a3fddc01080157fcc3ff36f5ca00ed;
mem[1020] = 144'h01cb008f008afdb2024a028502e3008f00a8;
mem[1021] = 144'h00fd011bfe370192018b00ecff55fe7a004b;
mem[1022] = 144'h05d805050088fe1effe700defd59fbe3fb10;
mem[1023] = 144'h00290102fec0007602beff0ffeb7fee8fad7;
end

always @ (posedge clk) begin
	q_a <= mem[addr_a];
end

always @ (posedge clk) begin
	q_b <= mem[addr_b];
end

endmodule