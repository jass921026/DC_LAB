`timescale 1ns/1ns

module wt_mem0 #(parameter ADDR_WIDTH = 11, DATA_WIDTH = 144, DEPTH = 76) (
input wire clk,
input wire [ADDR_WIDTH-1:0] addr_a, 
input wire [ADDR_WIDTH-1:0] addr_b, 
output reg [DATA_WIDTH-1:0] q_a,
output reg [DATA_WIDTH-1:0] q_b
);

reg [DATA_WIDTH-1:0] mem [0:DEPTH-1];

initial begin
mem[0] = 144'hfd180378f965f790f29519cc167f161107d0;
mem[1] = 144'h012c0bc122131042235b1f9bf3fbfaa60e2a;
mem[2] = 144'h0c170c9b0651ff180568fe90efd7f954f9d0;
mem[3] = 144'hfacafecbeef30cfa093f00ad08fd0b410860;
mem[4] = 144'h0b2d04e60616fe00fbb1fac5f701f651efd4;
mem[5] = 144'h07ed0237fea70df306b602d701a4039bfcb6;
mem[6] = 144'h045004dc082306580227fdb1f7d9fb34fd78;
mem[7] = 144'h00c3fb95f6450afb06b2044504bd03b00357;
mem[8] = 144'hf3faf9b000bb0fd60b3a06640d840144f898;
mem[9] = 144'hf244f3b1f789faccfda3011e0b960f030969;
mem[10] = 144'he7fffdb60965fa0f06a10f75113d13a702b4;
mem[11] = 144'hef89f82f009cf55103670627fc4c0950110b;
mem[12] = 144'hf65ef1ddfa9c000c07870eeb0595110c1265;
mem[13] = 144'hf60ef6b3f5b5f570f5d3ff63038301b903b5;
mem[14] = 144'h048e0db60abc0b440c32057ff66af246f57a;
mem[15] = 144'hfd9af71cf78e072201aa008b042409fa0441;
mem[16] = 144'hea8efc760057fc5e044cfcf500c5f56cef7d;
mem[17] = 144'h000d03c2116bf66707c312a5fd90ffb90519;
mem[18] = 144'h0142040e002c0d9d04d8014fff30fca6f4f2;
mem[19] = 144'hf703f9b1efe10890ff48fb240b8d0dbdfe89;
mem[20] = 144'h06450b0e02440000096c0114efe5f943fdb9;
mem[21] = 144'hffe3f9afee1f0da00500fbc70aa008b1ffc3;
mem[22] = 144'h0355f0e3e7b7f69fef56ed70f98df71ef3f3;
mem[23] = 144'h07b3f6e4f2630277f10cef080c40f293f20e;
mem[24] = 144'hfe48040b02af02ebfc6ffd2b027002de0192;
mem[25] = 144'hffc3ff4801ff000cf995ff96fb6c04050000;
mem[26] = 144'hfc87fe29ff7e0c5f0c66083b0bfc0428fd52;
mem[27] = 144'hf5f3f095f08bfd64016dfe1b0db40c5a0e37;
mem[28] = 144'hfe84fdb2ffa20c240ada0352023ff6fef72d;
mem[29] = 144'hfa6efbb9fe88fe56018dfe330a8302bf04eb;
mem[30] = 144'hf584f55ffd6204c50780071b0d2b10260d3a;
mem[31] = 144'hf3bbf55efc10f2dcf7ed045dfb72020e09ae;
mem[32] = 144'h0024033400b0fe2e001af7b7f084f606fc47;
mem[33] = 144'h06cbfd24fe8b060e087404a2091dfed1fb05;
mem[34] = 144'h064406240cea0432004a0389fb00fc13f8c5;
mem[35] = 144'hfe9bfc15fb6607e1102f060e055a0ab901ca;
mem[36] = 144'h0059fffa042306640f050c1208dc0b990a52;
mem[37] = 144'hf921fc5ff3060171040e003507670cdb0711;
mem[38] = 144'h05b00239060cf9d2fe3b0312ee91f370f099;
mem[39] = 144'h0784f6d6f58d11f10739fefd0425074105b7;
mem[40] = 144'h05110a5700730ce40e0d03a303ac031efbf3;
mem[41] = 144'hf79af9f8f0c106a3fe66fda012310c71023d;
mem[42] = 144'h069605b8034806230af600cffb2ff9aafa56;
mem[43] = 144'hfd3ff227f23f067304caf84a0781052a046e;
mem[44] = 144'hff01f7c8edb9f9cdf397f37701e3f81b00f4;
mem[45] = 144'h062101daf8a403defb82f6ba082ef580f7aa;
mem[46] = 144'hebebf7bf0144f119f951fc04f00000cdff7c;
mem[47] = 144'hf027055b11aced390b6d1372f88f0d770b76;
mem[48] = 144'h021bf71af145f8eaf179eff4f6edf701f3fd;
mem[49] = 144'h076ef490f54605c3fbd7ec020dc60015f847;
mem[50] = 144'hfa8bfe4602d1fc57032c0123ff3400c8fc72;
mem[51] = 144'h02240059012dfeed0069034a0002f9f9fc12;
mem[52] = 144'hef35fc4d01b4edeefc270640f92106c7093d;
mem[53] = 144'hfc4801980d25f31c087f08b1f15e0a720662;
mem[54] = 144'h005303c7fd7b0530030d0473fd500057ffc9;
mem[55] = 144'hfbda00c802af0024fe6cfddcfc2903ddfd00;
mem[56] = 144'h0b6304300e17e855eb88f89deccaf238f27e;
mem[57] = 144'h0c4b15cf1a1a0c8e09c9113ee731ed27f164;
mem[58] = 144'h08140b26035bfc56f79dfdace23fedcffada;
mem[59] = 144'h0c22061afa8013820a4e06dbf601fbebfa8f;
mem[60] = 144'hf722fdbefef8081b04e002f702c0fbf4fb41;
mem[61] = 144'hf893feff0209f970003ffce40f5e06a703bd;
mem[62] = 144'h0602ff80fee4fc8002f4fb2ff765f915fca1;
mem[63] = 144'hfb2000def5f207890526f92108fd0109fd43;
mem[64] = 144'h04670551ffb5016e0811ff5801b0f6b3f716;
mem[65] = 144'hfc98f7f0f72003c20736ff3c0adb0ad1fc90;
mem[66] = 144'h0456064dff92041c0670fce20a8d072bfa5b;
mem[67] = 144'h0404079dfb5e00a3fb23fc1efdaffcccfc4c;
mem[68] = 144'h09790312fb4300daff9303c207cb0023f2fc;
mem[69] = 144'h04f9f825fe46059ff712f978fa67fd2f00f6;
mem[70] = 144'hfbe7fc04fba60145082dfb35fdf4fd950690;
mem[71] = 144'hf4cbfebb06a2fb4ffec1fcde080ffd780172;
mem[72] = 144'h060d05adf8150639f49b0775066cfec2ff3b;
mem[73] = 144'hfc4b04ddfaae04910264fc29f18b00af08dc;
mem[74] = 144'h00400642fd0f01b802dbfc8a057801fd05a8;
mem[75] = 144'h0485fd59045bf9d505fcffccf78efe8bff14;
end

always @ (posedge clk) begin
	q_a <= mem[addr_a];
end

always @ (posedge clk) begin
	q_b <= mem[addr_b];
end

endmodule