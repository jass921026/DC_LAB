
module altpll (
	clk_clk,
	reset_reset_n,
	altpll_25m_clk_clk);	

	input		clk_clk;
	input		reset_reset_n;
	output		altpll_25m_clk_clk;
endmodule
