// Module for mouse communication

module Mouse
(
    input clk,  // system clock
    input rst,  // system reset
    inout ps2_clk,  // mouse clock
    inout ps2_data, // mouse data
    output [7:0] data,  // module output 
);

// Todo: Send reset, Send enable streaming, receive streaming input

endmodule