`timescale 1ns/1ns

module wt_mem3 #(parameter ADDR_WIDTH = 11, DATA_WIDTH = 144, DEPTH = 76) (
input wire clk,
input wire [ADDR_WIDTH-1:0] addr_a, 
input wire [ADDR_WIDTH-1:0] addr_b, 
output reg [DATA_WIDTH-1:0] q_a,
output reg [DATA_WIDTH-1:0] q_b
);

reg [DATA_WIDTH-1:0] mem [0:DEPTH-1];

initial begin
mem[0] = 144'h177b1829fd8016ec1cf4fe04167a1ed7f9b2;
mem[1] = 144'hf5c508f804ba04be170a1e740b9417640e0c;
mem[2] = 144'h03ec095bffb0095102c70974fcf5ffe306ec;
mem[3] = 144'h0a5a02fa03d509ca0ab60255fe2905bd029a;
mem[4] = 144'h071a08b505f703ed063cffe4faa5007505a6;
mem[5] = 144'h02b8048d0795019a08460560023103b000de;
mem[6] = 144'h0250043cfd430565071a0774049303a60594;
mem[7] = 144'h0648087dff2a072903a5ff86fdc405cf02ac;
mem[8] = 144'hfb4af496f7dbfa4f01a30588015004b50876;
mem[9] = 144'hf788f918fe8aff10082f02d0090909380092;
mem[10] = 144'hf766fbb9fcd7f35cfd5707d7fe4a0a280584;
mem[11] = 144'heeeff7f4018ff64506930aa3019b0b210bb0;
mem[12] = 144'h01ebf7a9f4dffd2bfab1fcde03a304df0b01;
mem[13] = 144'hf4d1fa44f2a0fa3bfe35059e01110d080b56;
mem[14] = 144'hf659f96a023207010233031f0258015b0098;
mem[15] = 144'h04a20888027f041b0b5f096903f804cafa59;
mem[16] = 144'hf56ffa57096ff2fe018e0315f97f01ff051c;
mem[17] = 144'hf272005e0c86f49b0685060d062d014a03ae;
mem[18] = 144'hfb5f049400060252048503de07bf03b405e1;
mem[19] = 144'h03b8043efb8908f7060afe2c07600217fce9;
mem[20] = 144'h0204feaaf811082d04890704fe0107ac06f2;
mem[21] = 144'h0317ff70fc2101b208210073fe8403a8f997;
mem[22] = 144'h026c082bf54b0b2908a6f59d046205fff33a;
mem[23] = 144'h0ab7f905f29d0608fab7ee16042ffbd7f4c2;
mem[24] = 144'hfce5fa77fee3fb1efe45fb650307fb99f987;
mem[25] = 144'hfb25ff01fa4dfee2fd4efbd8fb15fde9fdc4;
mem[26] = 144'hfa67f807f4f30601fc7a06680bbd09cc03c6;
mem[27] = 144'hf55ff398fb9a00bc02cf04ba04df0a1505bc;
mem[28] = 144'hf3aaff070326fd9608a4003bfe2902c40038;
mem[29] = 144'hfdb1042906f10002060505b108a90205ffff;
mem[30] = 144'hf782f212f72bfa8df921ffcc02770624039a;
mem[31] = 144'hf7c6f13efd7bf920fcd30261063707490e13;
mem[32] = 144'h06e90031028f0852025503ec040507e200f7;
mem[33] = 144'h05e5fe6a01760508023bfd7e0316f80af559;
mem[34] = 144'hfe6103e80549062901b5041dfde4005f049d;
mem[35] = 144'h068a05b7fff4014d082902e7007000adfd1f;
mem[36] = 144'h02e7ff4cfcd2027702ae0417ffef027f0b44;
mem[37] = 144'hfcc5fa3cff1105aa09db04f404500b240ab8;
mem[38] = 144'h0895ff0efa72028e081c04c0fbcb00370818;
mem[39] = 144'h0792011df8af0b0f0b3a002afc12fe6eff78;
mem[40] = 144'h0042fdf5fcbf03b106b006e8070801dd031c;
mem[41] = 144'h05bb035dfdb402b90817088605540758ffa8;
mem[42] = 144'hfdf70040f91c05400089085104c1064f0126;
mem[43] = 144'hfea500dafebf00d20744059c0210057a0539;
mem[44] = 144'h095903affd4907520003f507086401c1f471;
mem[45] = 144'h0258feaffbabfc62f488f5310322fa44f6c9;
mem[46] = 144'hfa61f5be083af3d8f8e1091bf447f758065a;
mem[47] = 144'hf81dfe400f94f29b04480e47f3cb06db04c9;
mem[48] = 144'h0ceb019cf6920c460418f2bd07690807f528;
mem[49] = 144'h0711f94ff92e08f4fd08f95e009001e4f5c3;
mem[50] = 144'hfd1d01d7fd2efd42fc0cfd8801d7fdf200c0;
mem[51] = 144'h022bfcd00078ff27fe77ff58fa77fead0312;
mem[52] = 144'hf989f9740523f426f5a3011af394f7d20c18;
mem[53] = 144'hf5d5fb350b1bf331ff2d0bcafae002cf0de9;
mem[54] = 144'h02a9faa702ed0166fb59fe45fb78fe7800db;
mem[55] = 144'hfea00445fab9ff95ffeb003800a5034a0247;
mem[56] = 144'h0be10db00904071afc2301edf415ee87f0ac;
mem[57] = 144'h081e0dbb0a7ffe22f70dfcd7eec6f275f1f8;
mem[58] = 144'h03b90b610a46feed00bd05fefe88fa64f913;
mem[59] = 144'h0af604d80788fee00a45ff82f103f25bf8e8;
mem[60] = 144'hf38dff550317fcc8043c03f4ffc509b706e6;
mem[61] = 144'hf527fdff074b024a021f05a0040502f500e7;
mem[62] = 144'h0489072c06b5ffe70a74012e053e021005b7;
mem[63] = 144'h0851052dfeb100ff08160215012d03ef044a;
mem[64] = 144'hfee9fe78fdfc05bb07ed09600603ff32ff51;
mem[65] = 144'h074c050701f806ae031201a1049203bffe40;
mem[66] = 144'hf968f86ffb8bff8f0204fd66f81cfc1203e0;
mem[67] = 144'hfdcbf81af8810a3b00e80734021bfa16fd59;
mem[68] = 144'h053eff65085004f8f95e077df9edfdd4fa23;
mem[69] = 144'h013d001af960fb16fac6f8a5fee600880b80;
mem[70] = 144'h075bf94ef62cfcc605faf344fc87f8b7f40a;
mem[71] = 144'hfab1fa50f2a0f49902aaf0f308a700d3016d;
mem[72] = 144'h01e2ff090491fddfffcdf8dcf2f9f82af253;
mem[73] = 144'hf8c5fc95083c0576fa650924fe28050ffe01;
mem[74] = 144'h067b069b0244019af8770586073b06070076;
mem[75] = 144'h038efbf0fc0afb67fcca046505a403d002a5;
end

always @ (posedge clk) begin
	q_a <= mem[addr_a];
end

always @ (posedge clk) begin
	q_b <= mem[addr_b];
end

endmodule