module generate_problem(
	input[7:0] problem_index,
	output[23:0] problem
);
	always_comb begin
		case(problem_index)
			8'd000:problem = 24'b111100011011000110100010;
			8'd001:problem = 24'b111100011100000110100000;
			8'd002:problem = 24'b111100011101000110100001;
			8'd003:problem = 24'b111100011110000110100001;
			8'd004:problem = 24'b111100011011001010100011;
			8'd005:problem = 24'b111100011101001010100010;
			8'd006:problem = 24'b111100011011001110100100;
			8'd007:problem = 24'b111100011101001110100011;
			8'd008:problem = 24'b111100011011010010100101;
			8'd009:problem = 24'b111100011101010010100100;
			8'd010:problem = 24'b111100011011010110100110;
			8'd011:problem = 24'b111100011101010110100101;
			8'd012:problem = 24'b111100011011011010100111;
			8'd013:problem = 24'b111100011101011010100110;
			8'd014:problem = 24'b111100011011011110101000;
			8'd015:problem = 24'b111100011101011110100111;
			8'd016:problem = 24'b111100011011100010101001;
			8'd017:problem = 24'b111100011101100010101000;
			8'd018:problem = 24'b111100011101100110101001;
			8'd019:problem = 24'b111100101011000110100011;
			8'd020:problem = 24'b111100101100000110100001;
			8'd021:problem = 24'b111100101101000110100010;
			8'd022:problem = 24'b111100101110000110100010;
			8'd023:problem = 24'b111100101011001010100100;
			8'd024:problem = 24'b111100101100001010100000;
			8'd025:problem = 24'b111100101101001010100100;
			8'd026:problem = 24'b111100101110001010100001;
			8'd027:problem = 24'b111100101011001110100101;
			8'd028:problem = 24'b111100101101001110100110;
			8'd029:problem = 24'b111100101011010010100110;
			8'd030:problem = 24'b111100101101010010101000;
			8'd031:problem = 24'b111100101011010110100111;
			8'd032:problem = 24'b111100101011011010101000;
			8'd033:problem = 24'b111100101011011110101001;
			8'd034:problem = 24'b111100111011000110100100;
			8'd035:problem = 24'b111100111100000110100010;
			8'd036:problem = 24'b111100111101000110100011;
			8'd037:problem = 24'b111100111110000110100011;
			8'd038:problem = 24'b111100111011001010100101;
			8'd039:problem = 24'b111100111100001010100001;
			8'd040:problem = 24'b111100111101001010100110;
			8'd041:problem = 24'b111100111011001110100110;
			8'd042:problem = 24'b111100111100001110100000;
			8'd043:problem = 24'b111100111101001110101001;
			8'd044:problem = 24'b111100111110001110100001;
			8'd045:problem = 24'b111100111011010010100111;
			8'd046:problem = 24'b111100111011010110101000;
			8'd047:problem = 24'b111100111011011010101001;
			8'd048:problem = 24'b111101001011000110100101;
			8'd049:problem = 24'b111101001100000110100011;
			8'd050:problem = 24'b111101001101000110100100;
			8'd051:problem = 24'b111101001110000110100100;
			8'd052:problem = 24'b111101001011001010100110;
			8'd053:problem = 24'b111101001100001010100010;
			8'd054:problem = 24'b111101001101001010101000;
			8'd055:problem = 24'b111101001110001010100010;
			8'd056:problem = 24'b111101001011001110100111;
			8'd057:problem = 24'b111101001100001110100001;
			8'd058:problem = 24'b111101001011010010101000;
			8'd059:problem = 24'b111101001100010010100000;
			8'd060:problem = 24'b111101001110010010100001;
			8'd061:problem = 24'b111101001011010110101001;
			8'd062:problem = 24'b111101011011000110100110;
			8'd063:problem = 24'b111101011100000110100100;
			8'd064:problem = 24'b111101011101000110100101;
			8'd065:problem = 24'b111101011110000110100101;
			8'd066:problem = 24'b111101011011001010100111;
			8'd067:problem = 24'b111101011100001010100011;
			8'd068:problem = 24'b111101011011001110101000;
			8'd069:problem = 24'b111101011100001110100010;
			8'd070:problem = 24'b111101011011010010101001;
			8'd071:problem = 24'b111101011100010010100001;
			8'd072:problem = 24'b111101011100010110100000;
			8'd073:problem = 24'b111101011110010110100001;
			8'd074:problem = 24'b111101101011000110100111;
			8'd075:problem = 24'b111101101100000110100101;
			8'd076:problem = 24'b111101101101000110100110;
			8'd077:problem = 24'b111101101110000110100110;
			8'd078:problem = 24'b111101101011001010101000;
			8'd079:problem = 24'b111101101100001010100100;
			8'd080:problem = 24'b111101101110001010100011;
			8'd081:problem = 24'b111101101011001110101001;
			8'd082:problem = 24'b111101101100001110100011;
			8'd083:problem = 24'b111101101110001110100010;
			8'd084:problem = 24'b111101101100010010100010;
			8'd085:problem = 24'b111101101100010110100001;
			8'd086:problem = 24'b111101101100011010100000;
			8'd087:problem = 24'b111101101110011010100001;
			8'd088:problem = 24'b111101111011000110101000;
			8'd089:problem = 24'b111101111100000110100110;
			8'd090:problem = 24'b111101111101000110100111;
			8'd091:problem = 24'b111101111110000110100111;
			8'd092:problem = 24'b111101111011001010101001;
			8'd093:problem = 24'b111101111100001010100101;
			8'd094:problem = 24'b111101111100001110100100;
			8'd095:problem = 24'b111101111100010010100011;
			8'd096:problem = 24'b111101111100010110100010;
			8'd097:problem = 24'b111101111100011010100001;
			8'd098:problem = 24'b111101111100011110100000;
			8'd099:problem = 24'b111101111110011110100001;
			8'd100:problem = 24'b111110001011000110101001;
			8'd101:problem = 24'b111110001100000110100111;
			8'd102:problem = 24'b111110001101000110101000;
			8'd103:problem = 24'b111110001110000110101000;
			8'd104:problem = 24'b111110001100001010100110;
			8'd105:problem = 24'b111110001110001010100100;
			8'd106:problem = 24'b111110001100001110100101;
			8'd107:problem = 24'b111110001100010010100100;
			8'd108:problem = 24'b111110001110010010100010;
			8'd109:problem = 24'b111110001100010110100011;
			8'd110:problem = 24'b111110001100011010100010;
			8'd111:problem = 24'b111110001100011110100001;
			8'd112:problem = 24'b111110001100100010100000;
			8'd113:problem = 24'b111110001110100010100001;
			8'd114:problem = 24'b111110011100000110101000;
			8'd115:problem = 24'b111110011101000110101001;
			8'd116:problem = 24'b111110011110000110101001;
			8'd117:problem = 24'b111110011100001010100111;
			8'd118:problem = 24'b111110011100001110100110;
			8'd119:problem = 24'b111110011110001110100011;
			8'd120:problem = 24'b111110011100010010100101;
			8'd121:problem = 24'b111110011100010110100100;
			8'd122:problem = 24'b111110011100011010100011;
			8'd123:problem = 24'b111110011100011110100010;
			8'd124:problem = 24'b111110011100100010100001;
			8'd125:problem = 24'b111110011100100110100000;
			8'd126:problem = 24'b111110011110100110100001;
			8'd127:problem = 24'b000100001100000110101001;
			8'd128:problem = 24'b000100001100001010101000;
			8'd129:problem = 24'b000100001110001010100101;
			8'd130:problem = 24'b000100001100001110100111;
			8'd131:problem = 24'b000100001100010010100110;
			8'd132:problem = 24'b000100001100010110100101;
			8'd133:problem = 24'b000100001110010110100010;
			8'd134:problem = 24'b000100001100011010100100;
			8'd135:problem = 24'b000100001100011110100011;
			8'd136:problem = 24'b000100001100100010100010;
			8'd137:problem = 24'b000100001100100110100001;
			8'd138:problem = 24'b000100011100001010101001;
			8'd139:problem = 24'b000100011100001110101000;
			8'd140:problem = 24'b000100011100010010100111;
			8'd141:problem = 24'b000100011100010110100110;
			8'd142:problem = 24'b000100011100011010100101;
			8'd143:problem = 24'b000100011100011110100100;
			8'd144:problem = 24'b000100011100100010100011;
			8'd145:problem = 24'b000100011100100110100010;
			8'd146:problem = 24'b000100101110001010100110;
			8'd147:problem = 24'b000100101100001110101001;
			8'd148:problem = 24'b000100101110001110100100;
			8'd149:problem = 24'b000100101100010010101000;
			8'd150:problem = 24'b000100101110010010100011;
			8'd151:problem = 24'b000100101100010110100111;
			8'd152:problem = 24'b000100101100011010100110;
			8'd153:problem = 24'b000100101110011010100010;
			8'd154:problem = 24'b000100101100011110100101;
			8'd155:problem = 24'b000100101100100010100100;
			8'd156:problem = 24'b000100101100100110100011;
			8'd157:problem = 24'b000100111100010010101001;
			8'd158:problem = 24'b000100111100010110101000;
			8'd159:problem = 24'b000100111100011010100111;
			8'd160:problem = 24'b000100111100011110100110;
			8'd161:problem = 24'b000100111100100010100101;
			8'd162:problem = 24'b000100111100100110100100;
			8'd163:problem = 24'b000101001110001010100111;
			8'd164:problem = 24'b000101001100010110101001;
			8'd165:problem = 24'b000101001100011010101000;
			8'd166:problem = 24'b000101001100011110100111;
			8'd167:problem = 24'b000101001110011110100010;
			8'd168:problem = 24'b000101001100100010100110;
			8'd169:problem = 24'b000101001100100110100101;
			8'd170:problem = 24'b000101011110001110100101;
			8'd171:problem = 24'b000101011110010110100011;
			8'd172:problem = 24'b000101011100011010101001;
			8'd173:problem = 24'b000101011100011110101000;
			8'd174:problem = 24'b000101011100100010100111;
			8'd175:problem = 24'b000101011100100110100110;
			8'd176:problem = 24'b000101101110001010101000;
			8'd177:problem = 24'b000101101110010010100100;
			8'd178:problem = 24'b000101101100011110101001;
			8'd179:problem = 24'b000101101100100010101000;
			8'd180:problem = 24'b000101101110100010100010;
			8'd181:problem = 24'b000101101100100110100111;
			8'd182:problem = 24'b000101111100100010101001;
			8'd183:problem = 24'b000101111100100110101000;
			8'd184:problem = 24'b000110001110001010101001;
			8'd185:problem = 24'b000110001110001110100110;
			8'd186:problem = 24'b000110001110011010100011;
			8'd187:problem = 24'b000110001100100110101001;
			8'd188:problem = 24'b000110001110100110100010;
			8'd189:problem = 24'b001000001110010010100101;
			8'd190:problem = 24'b001000001110010110100100;
			8'd191:problem = 24'b001000011110001110100111;
			8'd192:problem = 24'b001000011110011110100011;
			8'd193:problem = 24'b001001001110001110101000;
			8'd194:problem = 24'b001001001110010010100110;
			8'd195:problem = 24'b001001001110011010100100;
			8'd196:problem = 24'b001001001110100010100011;
			8'd197:problem = 24'b001001011110010110100101;
			8'd198:problem = 24'b001001111110001110101001;
			8'd199:problem = 24'b001001111110100110100011;
			8'd200:problem = 24'b001010001110010010100111;
			8'd201:problem = 24'b001010001110011110100100;
			8'd202:problem = 24'b001100001110010110100110;
			8'd203:problem = 24'b001100001110011010100101;
			8'd204:problem = 24'b001100101110010010101000;
			8'd205:problem = 24'b001100101110100010100100;
			8'd206:problem = 24'b001101011110010110100111;
			8'd207:problem = 24'b001101011110011110100101;
			8'd208:problem = 24'b001101101110010010101001;
			8'd209:problem = 24'b001101101110011010100110;
			8'd210:problem = 24'b001101101110100110100100;
			8'd211:problem = 24'b010000001110010110101000;
			8'd212:problem = 24'b010000001110100010100101;
			8'd213:problem = 24'b010000101110011010100111;
			8'd214:problem = 24'b010000101110011110100110;
			8'd215:problem = 24'b010001011110010110101001;
			8'd216:problem = 24'b010001011110100110100101;
			8'd217:problem = 24'b010010001110011010101000;
			8'd218:problem = 24'b010010001110100010100110;
			8'd219:problem = 24'b010010011110011110100111;
			8'd220:problem = 24'b010101001110011010101001;
			8'd221:problem = 24'b010101001110100110100110;
			8'd222:problem = 24'b010101101110011110101000;
			8'd223:problem = 24'b010101101110100010100111;
			8'd224:problem = 24'b011000111110011110101001;
			8'd225:problem = 24'b011000111110100110100111;
			8'd226:problem = 24'b011001001110100010101000;
			8'd227:problem = 24'b011100101110100010101001;
			8'd228:problem = 24'b011100101110100110101000;
			default:problem = 24'b0;
		endcase
	end
endmodule
